// Copyright 2022 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Fabian Schuiki <fschuiki@iis.ee.ethz.ch>
// Florian Zaruba <zarubaf@iis.ee.ethz.ch>
// Stefan Mach <smach@iis.ee.ethz.ch>
// Thomas Benz <tbenz@iis.ee.ethz.ch>
// Paul Scheffler <paulsc@iis.ee.ethz.ch>
// Wolfgang Roenninger <wroennin@iis.ee.ethz.ch>
//
// AUTOMATICALLY GENERATED by gen_bootrom.py; edit the script instead.

module cheshire_bootrom #(
    parameter int unsigned AddrWidth = 32,
    parameter int unsigned DataWidth = 32
)(
    input  logic                 clk_i,
    input  logic                 rst_ni,
    input  logic                 req_i,
    input  logic [AddrWidth-1:0] addr_i,
    output logic [DataWidth-1:0] data_o
);
    localparam unsigned NumWords = 2048;
    logic [$clog2(NumWords)-1:0] word;

    assign word = addr_i / (DataWidth / 8);

    always_comb begin
        data_o = '0;
        unique case (word)
        000: data_o = 32'h42014081 /* 0x0000 */;
            001: data_o = 32'h43014281 /* 0x0004 */;
            002: data_o = 32'h44014381 /* 0x0008 */;
            003: data_o = 32'h45014481 /* 0x000c */;
            004: data_o = 32'h46014581 /* 0x0010 */;
            005: data_o = 32'h47014681 /* 0x0014 */;
            006: data_o = 32'h48014781 /* 0x0018 */;
            007: data_o = 32'h49014881 /* 0x001c */;
            008: data_o = 32'h4a014981 /* 0x0020 */;
            009: data_o = 32'h4b014a81 /* 0x0024 */;
            010: data_o = 32'h4c014b81 /* 0x0028 */;
            011: data_o = 32'h4d014c81 /* 0x002c */;
            012: data_o = 32'h4e014d81 /* 0x0030 */;
            013: data_o = 32'h4f014e81 /* 0x0034 */;
            014: data_o = 32'h43214f81 /* 0x0038 */;
            015: data_o = 32'h30431073 /* 0x003c */;
            016: data_o = 32'h23734281 /* 0x0040 */;
            017: data_o = 32'h9663f140 /* 0x0044 */;
            018: data_o = 32'h01170a62 /* 0x0048 */;
            019: data_o = 32'h01130e01 /* 0x004c */;
            020: data_o = 32'h2197fae1 /* 0x0050 */;
            021: data_o = 32'h81930000 /* 0x0054 */;
            022: data_o = 32'h0297bc21 /* 0x0058 */;
            023: data_o = 32'h82930100 /* 0x005c */;
            024: data_o = 32'ha283fa62 /* 0x0060 */;
            025: data_o = 32'hf2930502 /* 0x0064 */;
            026: data_o = 32'h8e630022 /* 0x0068 */;
            027: data_o = 32'h12970202 /* 0x006c */;
            028: data_o = 32'h82930100 /* 0x0070 */;
            029: data_o = 32'ha303f922 /* 0x0074 */;
            030: data_o = 32'h0ee30482 /* 0x0078 */;
            031: data_o = 32'h537dfe03 /* 0x007c */;
            032: data_o = 32'h0062a023 /* 0x0080 */;
            033: data_o = 32'h0062a223 /* 0x0084 */;
            034: data_o = 32'ha8234305 /* 0x0088 */;
            035: data_o = 32'h02970062 /* 0x008c */;
            036: data_o = 32'h82930100 /* 0x0090 */;
            037: data_o = 32'h0117f722 /* 0x0094 */;
            038: data_o = 32'h01130e00 /* 0x0098 */;
            039: data_o = 32'ha283f6a1 /* 0x009c */;
            040: data_o = 32'h91160542 /* 0x00a0 */;
            041: data_o = 32'h02971161 /* 0x00a4 */;
            042: data_o = 32'h82930100 /* 0x00a8 */;
            043: data_o = 32'ha283f5a2 /* 0x00ac */;
            044: data_o = 32'h81630482 /* 0x00b0 */;
            045: data_o = 32'h92820a02 /* 0x00b4 */;
            046: data_o = 32'h01000297 /* 0x00b8 */;
            047: data_o = 32'hf4828293 /* 0x00bc */;
            048: data_o = 32'h00a2a823 /* 0x00c0 */;
            049: data_o = 32'haa239101 /* 0x00c4 */;
            050: data_o = 32'h000f00a2 /* 0x00c8 */;
            051: data_o = 32'h02970ff0 /* 0x00cc */;
            052: data_o = 32'h82930004 /* 0x00d0 */;
            053: data_o = 32'h0397f322 /* 0x00d4 */;
            054: data_o = 32'h83930100 /* 0x00d8 */;
            055: data_o = 32'ha383f2a3 /* 0x00dc */;
            056: data_o = 32'h038a04c3 /* 0x00e0 */;
            057: data_o = 32'h43059396 /* 0x00e4 */;
            058: data_o = 32'h0062a023 /* 0x00e8 */;
            059: data_o = 32'hcce30291 /* 0x00ec */;
            060: data_o = 32'h0073fe72 /* 0x00f0 */;
            061: data_o = 32'h23731050 /* 0x00f4 */;
            062: data_o = 32'h73133440 /* 0x00f8 */;
            063: data_o = 32'h0ae30083 /* 0x00fc */;
            064: data_o = 32'h0297fe03 /* 0x0100 */;
            065: data_o = 32'h82930004 /* 0x0104 */;
            066: data_o = 32'h2373efe2 /* 0x0108 */;
            067: data_o = 32'h030af140 /* 0x010c */;
            068: data_o = 32'h20239316 /* 0x0110 */;
            069: data_o = 32'h03970003 /* 0x0114 */;
            070: data_o = 32'h83930100 /* 0x0118 */;
            071: data_o = 32'ha383eea3 /* 0x011c */;
            072: data_o = 32'h038a04c3 /* 0x0120 */;
            073: data_o = 32'ha3039396 /* 0x0124 */;
            074: data_o = 32'h1ee30002 /* 0x0128 */;
            075: data_o = 32'h0291fe03 /* 0x012c */;
            076: data_o = 32'hfe72cbe3 /* 0x0130 */;
            077: data_o = 32'h01000297 /* 0x0134 */;
            078: data_o = 32'hecc28293 /* 0x0138 */;
            079: data_o = 32'h0142e303 /* 0x013c */;
            080: data_o = 32'he2831302 /* 0x0140 */;
            081: data_o = 32'he2b30102 /* 0x0144 */;
            082: data_o = 32'h25730062 /* 0x0148 */;
            083: data_o = 32'h80e7f140 /* 0x014c */;
            084: data_o = 32'h80820002 /* 0x0150 */;
            085: data_o = 32'h43014281 /* 0x0154 */;
            086: data_o = 32'h0ff0000f /* 0x0158 */;
            087: data_o = 32'h0000100f /* 0x015c */;
            088: data_o = 32'h031010ef /* 0x0160 */;
            089: data_o = 32'h65130506 /* 0x0164 */;
            090: data_o = 32'h02970015 /* 0x0168 */;
            091: data_o = 32'h82930100 /* 0x016c */;
            092: data_o = 32'ha423e962 /* 0x0170 */;
            093: data_o = 32'h900200a2 /* 0x0174 */;
            094: data_o = 32'h10500073 /* 0x0178 */;
            095: data_o = 32'h171bbff5 /* 0x017c */;
            096: data_o = 32'h579b0185 /* 0x0180 */;
            097: data_o = 32'h66c10185 /* 0x0184 */;
            098: data_o = 32'h86938fd9 /* 0x0188 */;
            099: data_o = 32'h571bf006 /* 0x018c */;
            100: data_o = 32'h8f750085 /* 0x0190 */;
            101: data_o = 32'h151b8fd9 /* 0x0194 */;
            102: data_o = 32'h07370085 /* 0x0198 */;
            103: data_o = 32'h8d7900ff /* 0x019c */;
            104: data_o = 32'h80828d5d /* 0x01a0 */;
            105: data_o = 32'hc611832a /* 0x01a4 */;
            106: data_o = 32'h00b30023 /* 0x01a8 */;
            107: data_o = 32'h0305167d /* 0x01ac */;
            108: data_o = 32'h8082fe65 /* 0x01b0 */;
            109: data_o = 32'hca09832a /* 0x01b4 */;
            110: data_o = 32'h00058383 /* 0x01b8 */;
            111: data_o = 32'h00730023 /* 0x01bc */;
            112: data_o = 32'h0305167d /* 0x01c0 */;
            113: data_o = 32'hfa6d0585 /* 0x01c4 */;
            114: data_o = 32'h0b638082 /* 0x01c8 */;
            115: data_o = 32'h87631605 /* 0x01cc */;
            116: data_o = 32'hd7b71605 /* 0x01d0 */;
            117: data_o = 32'h87933b9a /* 0x01d4 */;
            118: data_o = 32'hd5b3a007 /* 0x01d8 */;
            119: data_o = 32'h381702b7 /* 0x01dc */;
            120: data_o = 32'h08130100 /* 0x01e0 */;
            121: data_o = 32'h2303e228 /* 0x01e4 */;
            122: data_o = 32'h3e170108 /* 0x01e8 */;
            123: data_o = 32'h0e130100 /* 0x01ec */;
            124: data_o = 32'h3817e16e /* 0x01f0 */;
            125: data_o = 32'h30230100 /* 0x01f4 */;
            126: data_o = 32'h731301c5 /* 0x01f8 */;
            127: data_o = 32'h0813ffe3 /* 0x01fc */;
            128: data_o = 32'h3517e0e8 /* 0x0200 */;
            129: data_o = 32'h28230100 /* 0x0204 */;
            130: data_o = 32'h05130068 /* 0x0208 */;
            131: data_o = 32'h2303dfe5 /* 0x020c */;
            132: data_o = 32'h38170205 /* 0x0210 */;
            133: data_o = 32'h08130100 /* 0x0214 */;
            134: data_o = 32'h6313dee8 /* 0x0218 */;
            135: data_o = 32'h35170803 /* 0x021c */;
            136: data_o = 32'h20230100 /* 0x0220 */;
            137: data_o = 32'h05130268 /* 0x0224 */;
            138: data_o = 32'h2303de25 /* 0x0228 */;
            139: data_o = 32'h38170205 /* 0x022c */;
            140: data_o = 32'h08130100 /* 0x0230 */;
            141: data_o = 32'h6313dd28 /* 0x0234 */;
            142: data_o = 32'h35170023 /* 0x0238 */;
            143: data_o = 32'h20230100 /* 0x023c */;
            144: data_o = 32'h05130268 /* 0x0240 */;
            145: data_o = 32'h2303dc65 /* 0x0244 */;
            146: data_o = 32'h38170205 /* 0x0248 */;
            147: data_o = 32'h08130100 /* 0x024c */;
            148: data_o = 32'h6313db68 /* 0x0250 */;
            149: data_o = 32'h35170013 /* 0x0254 */;
            150: data_o = 32'h20230100 /* 0x0258 */;
            151: data_o = 32'h05130268 /* 0x025c */;
            152: data_o = 32'h2803daa5 /* 0x0260 */;
            153: data_o = 32'h67850205 /* 0x0264 */;
            154: data_o = 32'h01003517 /* 0x0268 */;
            155: data_o = 32'hd9850513 /* 0x026c */;
            156: data_o = 32'h10086813 /* 0x0270 */;
            157: data_o = 32'h51300893 /* 0x0274 */;
            158: data_o = 32'h9c37879b /* 0x0278 */;
            159: data_o = 32'h06300713 /* 0x027c */;
            160: data_o = 32'h03052023 /* 0x0280 */;
            161: data_o = 32'h12b00693 /* 0x0284 */;
            162: data_o = 32'h25700613 /* 0x0288 */;
            163: data_o = 32'h02b8d83b /* 0x028c */;
            164: data_o = 32'h02b7d7bb /* 0x0290 */;
            165: data_o = 32'h0018051b /* 0x0294 */;
            166: data_o = 32'h0105151b /* 0x0298 */;
            167: data_o = 32'h02b7573b /* 0x029c */;
            168: data_o = 32'h410787bb /* 0x02a0 */;
            169: data_o = 32'h02b6d6bb /* 0x02a4 */;
            170: data_o = 32'h9f990705 /* 0x02a8 */;
            171: data_o = 32'h02b6563b /* 0x02ac */;
            172: data_o = 32'h9f950685 /* 0x02b0 */;
            173: data_o = 32'h03079813 /* 0x02b4 */;
            174: data_o = 32'h03085813 /* 0x02b8 */;
            175: data_o = 32'h00160593 /* 0x02bc */;
            176: data_o = 32'h6b63862e /* 0x02c0 */;
            177: data_o = 32'h65c106b8 /* 0x02c4 */;
            178: data_o = 32'h25852601 /* 0x02c8 */;
            179: data_o = 32'h02b605bb /* 0x02cc */;
            180: data_o = 32'h93c117c2 /* 0x02d0 */;
            181: data_o = 32'h01003897 /* 0x02d4 */;
            182: data_o = 32'h27018fc9 /* 0x02d8 */;
            183: data_o = 32'hd2c88893 /* 0x02dc */;
            184: data_o = 32'h0106969b /* 0x02e0 */;
            185: data_o = 32'h01003817 /* 0x02e4 */;
            186: data_o = 32'h02f8a823 /* 0x02e8 */;
            187: data_o = 32'h08138ed9 /* 0x02ec */;
            188: data_o = 32'h3797d1c8 /* 0x02f0 */;
            189: data_o = 32'h2a230100 /* 0x02f4 */;
            190: data_o = 32'h879302d8 /* 0x02f8 */;
            191: data_o = 32'h6841d0e7 /* 0x02fc */;
            192: data_o = 32'h01003697 /* 0x0300 */;
            193: data_o = 32'h6733df8c /* 0x0304 */;
            194: data_o = 32'h86930107 /* 0x0308 */;
            195: data_o = 32'h3797d006 /* 0x030c */;
            196: data_o = 32'hded80100 /* 0x0310 */;
            197: data_o = 32'h87138d51 /* 0x0314 */;
            198: data_o = 32'h3797cf27 /* 0x0318 */;
            199: data_o = 32'hc3280100 /* 0x031c */;
            200: data_o = 32'hce678793 /* 0x0320 */;
            201: data_o = 32'h37974b98 /* 0x0324 */;
            202: data_o = 32'h87930100 /* 0x0328 */;
            203: data_o = 32'h6713cda7 /* 0x032c */;
            204: data_o = 32'hcb980017 /* 0x0330 */;
            205: data_o = 32'h80824501 /* 0x0334 */;
            206: data_o = 32'hb77187ae /* 0x0338 */;
            207: data_o = 32'h80824549 /* 0x033c */;
            208: data_o = 32'h80824545 /* 0x0340 */;
            209: data_o = 32'h07176631 /* 0x0344 */;
            210: data_o = 32'h07970004 /* 0x0348 */;
            211: data_o = 32'h07130004 /* 0x034c */;
            212: data_o = 32'h8793cba7 /* 0x0350 */;
            213: data_o = 32'h97b2cb67 /* 0x0354 */;
            214: data_o = 32'h27039732 /* 0x0358 */;
            215: data_o = 32'ha683ffc7 /* 0x035c */;
            216: data_o = 32'h1793ff87 /* 0x0360 */;
            217: data_o = 32'h97130207 /* 0x0364 */;
            218: data_o = 32'h93010206 /* 0x0368 */;
            219: data_o = 32'hece38fd9 /* 0x036c */;
            220: data_o = 32'h8082fca7 /* 0x0370 */;
            221: data_o = 32'hce85c929 /* 0x0374 */;
            222: data_o = 32'hffd6079b /* 0x0378 */;
            223: data_o = 32'h74634709 /* 0x037c */;
            224: data_o = 32'h076304f7 /* 0x0380 */;
            225: data_o = 32'h167d04e6 /* 0x0384 */;
            226: data_o = 32'h00c03633 /* 0x0388 */;
            227: data_o = 32'h25814781 /* 0x038c */;
            228: data_o = 32'h0086161b /* 0x0390 */;
            229: data_o = 32'h969b4701 /* 0x0394 */;
            230: data_o = 32'h979b00c6 /* 0x0398 */;
            231: data_o = 32'h8fd50097 /* 0x039c */;
            232: data_o = 32'h61188fd9 /* 0x03a0 */;
            233: data_o = 32'h8fcd8fd1 /* 0x03a4 */;
            234: data_o = 32'h4501cf5c /* 0x03a8 */;
            235: data_o = 32'h47898082 /* 0x03ac */;
            236: data_o = 32'h00f60d63 /* 0x03b0 */;
            237: data_o = 32'h18e3478d /* 0x03b4 */;
            238: data_o = 32'h2581fcf6 /* 0x03b8 */;
            239: data_o = 32'h46014781 /* 0x03bc */;
            240: data_o = 32'h40000713 /* 0x03c0 */;
            241: data_o = 32'h450dbfc9 /* 0x03c4 */;
            242: data_o = 32'h46018082 /* 0x03c8 */;
            243: data_o = 32'hb7c14785 /* 0x03cc */;
            244: data_o = 32'h46014785 /* 0x03d0 */;
            245: data_o = 32'h715dbf6d /* 0x03d4 */;
            246: data_o = 32'hf84afc26 /* 0x03d8 */;
            247: data_o = 32'hf052f44e /* 0x03dc */;
            248: data_o = 32'he486ec56 /* 0x03e0 */;
            249: data_o = 32'h892e84aa /* 0x03e4 */;
            250: data_o = 32'h89b68a32 /* 0x03e8 */;
            251: data_o = 32'he8918aba /* 0x03ec */;
            252: data_o = 32'h60a6450d /* 0x03f0 */;
            253: data_o = 32'h794274e2 /* 0x03f4 */;
            254: data_o = 32'h7a0279a2 /* 0x03f8 */;
            255: data_o = 32'h61616ae2 /* 0x03fc */;
            256: data_o = 32'he0a28082 /* 0x0400 */;
            257: data_o = 32'he85a6080 /* 0x0404 */;
            258: data_o = 32'he062e45e /* 0x0408 */;
            259: data_o = 32'hf813505c /* 0x040c */;
            260: data_o = 32'h278107f7 /* 0x0410 */;
            261: data_o = 32'hfe081ce3 /* 0x0414 */;
            262: data_o = 32'h0107d81b /* 0x0418 */;
            263: data_o = 32'h0087d89b /* 0x041c */;
            264: data_o = 32'h01186833 /* 0x0420 */;
            265: data_o = 32'h0187d79b /* 0x0424 */;
            266: data_o = 32'h00f867b3 /* 0x0428 */;
            267: data_o = 32'h07f7f793 /* 0x042c */;
            268: data_o = 32'h0717fff1 /* 0x0430 */;
            269: data_o = 32'h07970004 /* 0x0434 */;
            270: data_o = 32'h66310004 /* 0x0438 */;
            271: data_o = 32'hbce70713 /* 0x043c */;
            272: data_o = 32'hbca78793 /* 0x0440 */;
            273: data_o = 32'h97b29732 /* 0x0444 */;
            274: data_o = 32'hffc72583 /* 0x0448 */;
            275: data_o = 32'hff87a783 /* 0x044c */;
            276: data_o = 32'h17821582 /* 0x0450 */;
            277: data_o = 32'h8ddd9381 /* 0x0454 */;
            278: data_o = 32'h08170585 /* 0x0458 */;
            279: data_o = 32'h07970004 /* 0x045c */;
            280: data_o = 32'h08130004 /* 0x0460 */;
            281: data_o = 32'h8793ba68 /* 0x0464 */;
            282: data_o = 32'h97b2ba27 /* 0x0468 */;
            283: data_o = 32'h27039832 /* 0x046c */;
            284: data_o = 32'ha683ffc8 /* 0x0470 */;
            285: data_o = 32'h1793ff87 /* 0x0474 */;
            286: data_o = 32'h97130207 /* 0x0478 */;
            287: data_o = 32'h93010206 /* 0x047c */;
            288: data_o = 32'hece38fd9 /* 0x0480 */;
            289: data_o = 32'h481cfcb7 /* 0x0484 */;
            290: data_o = 32'h46014685 /* 0x0488 */;
            291: data_o = 32'hc81c9bf9 /* 0x048c */;
            292: data_o = 32'h0a000593 /* 0x0490 */;
            293: data_o = 32'hf0ef8526 /* 0x0494 */;
            294: data_o = 32'he125edff /* 0x0498 */;
            295: data_o = 32'h008a5593 /* 0x049c */;
            296: data_o = 32'hf5934685 /* 0x04a0 */;
            297: data_o = 32'h86360ff5 /* 0x04a4 */;
            298: data_o = 32'hf0ef8526 /* 0x04a8 */;
            299: data_o = 32'he531ecbf /* 0x04ac */;
            300: data_o = 32'h063b4609 /* 0x04b0 */;
            301: data_o = 32'h46854156 /* 0x04b4 */;
            302: data_o = 32'h0ffa7593 /* 0x04b8 */;
            303: data_o = 32'hf0ef8526 /* 0x04bc */;
            304: data_o = 32'hed05eb7f /* 0x04c0 */;
            305: data_o = 32'h040a8063 /* 0x04c4 */;
            306: data_o = 32'hfff98c13 /* 0x04c8 */;
            307: data_o = 32'h02000793 /* 0x04cc */;
            308: data_o = 32'hf3638be2 /* 0x04d0 */;
            309: data_o = 32'h8bbe0187 /* 0x04d4 */;
            310: data_o = 32'h0a0c0463 /* 0x04d8 */;
            311: data_o = 32'ha0194b01 /* 0x04dc */;
            312: data_o = 32'h077b7963 /* 0x04e0 */;
            313: data_o = 32'h016907b3 /* 0x04e4 */;
            314: data_o = 32'h0007c583 /* 0x04e8 */;
            315: data_o = 32'h86364685 /* 0x04ec */;
            316: data_o = 32'hf0ef8526 /* 0x04f0 */;
            317: data_o = 32'h0b05e83f /* 0x04f4 */;
            318: data_o = 32'h6406d565 /* 0x04f8 */;
            319: data_o = 32'h6ba26b42 /* 0x04fc */;
            320: data_o = 32'hb5fd6c02 /* 0x0500 */;
            321: data_o = 32'h46014685 /* 0x0504 */;
            322: data_o = 32'h0a100593 /* 0x0508 */;
            323: data_o = 32'hf0ef8526 /* 0x050c */;
            324: data_o = 32'hf565e67f /* 0x0510 */;
            325: data_o = 32'h460d4681 /* 0x0514 */;
            326: data_o = 32'h0ff9f593 /* 0x0518 */;
            327: data_o = 32'hf0ef8526 /* 0x051c */;
            328: data_o = 32'hfd61e57f /* 0x0520 */;
            329: data_o = 32'he793481c /* 0x0524 */;
            330: data_o = 32'hc81c0017 /* 0x0528 */;
            331: data_o = 32'hd79b505c /* 0x052c */;
            332: data_o = 32'hf7930107 /* 0x0530 */;
            333: data_o = 32'hebe307f7 /* 0x0534 */;
            334: data_o = 32'h99caff37 /* 0x0538 */;
            335: data_o = 32'h4f9c609c /* 0x053c */;
            336: data_o = 32'h04632781 /* 0x0540 */;
            337: data_o = 32'h00230009 /* 0x0544 */;
            338: data_o = 32'h090500f9 /* 0x0548 */;
            339: data_o = 32'hff2998e3 /* 0x054c */;
            340: data_o = 32'h9c4aa015 /* 0x0550 */;
            341: data_o = 32'h000c4583 /* 0x0554 */;
            342: data_o = 32'h86364685 /* 0x0558 */;
            343: data_o = 32'hf0ef8526 /* 0x055c */;
            344: data_o = 32'hfd41e17f /* 0x0560 */;
            345: data_o = 32'h0713481c /* 0x0564 */;
            346: data_o = 32'he7930200 /* 0x0568 */;
            347: data_o = 32'hc81c0017 /* 0x056c */;
            348: data_o = 32'h03376563 /* 0x0570 */;
            349: data_o = 32'h6b426406 /* 0x0574 */;
            350: data_o = 32'h6c026ba2 /* 0x0578 */;
            351: data_o = 32'hbd954501 /* 0x057c */;
            352: data_o = 32'h00094583 /* 0x0580 */;
            353: data_o = 32'h85264685 /* 0x0584 */;
            354: data_o = 32'hf0ef8636 /* 0x0588 */;
            355: data_o = 32'hf535debf /* 0x058c */;
            356: data_o = 32'he793481c /* 0x0590 */;
            357: data_o = 32'hc81c0017 /* 0x0594 */;
            358: data_o = 32'h994ebff1 /* 0x0598 */;
            359: data_o = 32'h64069a4e /* 0x059c */;
            360: data_o = 32'h6ba26b42 /* 0x05a0 */;
            361: data_o = 32'h19816c02 /* 0x05a4 */;
            362: data_o = 32'he40484e3 /* 0x05a8 */;
            363: data_o = 32'h7139bd99 /* 0x05ac */;
            364: data_o = 32'hf426f822 /* 0x05b0 */;
            365: data_o = 32'hec4ef04a /* 0x05b4 */;
            366: data_o = 32'hfc06e852 /* 0x05b8 */;
            367: data_o = 32'h03f67413 /* 0x05bc */;
            368: data_o = 32'h84b68932 /* 0x05c0 */;
            369: data_o = 32'h8a2e89aa /* 0x05c4 */;
            370: data_o = 32'he456ec31 /* 0x05c8 */;
            371: data_o = 32'h04000a93 /* 0x05cc */;
            372: data_o = 32'h00946563 /* 0x05d0 */;
            373: data_o = 32'h7d63a835 /* 0x05d4 */;
            374: data_o = 32'h86b30294 /* 0x05d8 */;
            375: data_o = 32'h47014084 /* 0x05dc */;
            376: data_o = 32'h00890633 /* 0x05e0 */;
            377: data_o = 32'h008a05b3 /* 0x05e4 */;
            378: data_o = 32'hf463854e /* 0x05e8 */;
            379: data_o = 32'h069300da /* 0x05ec */;
            380: data_o = 32'hf0ef0400 /* 0x05f0 */;
            381: data_o = 32'h0413de5f /* 0x05f4 */;
            382: data_o = 32'hdd710404 /* 0x05f8 */;
            383: data_o = 32'h70e26aa2 /* 0x05fc */;
            384: data_o = 32'h74a27442 /* 0x0600 */;
            385: data_o = 32'h69e27902 /* 0x0604 */;
            386: data_o = 32'h450d6a42 /* 0x0608 */;
            387: data_o = 32'h80826121 /* 0x060c */;
            388: data_o = 32'h744270e2 /* 0x0610 */;
            389: data_o = 32'h74a26aa2 /* 0x0614 */;
            390: data_o = 32'h69e27902 /* 0x0618 */;
            391: data_o = 32'h45016a42 /* 0x061c */;
            392: data_o = 32'h80826121 /* 0x0620 */;
            393: data_o = 32'h04000793 /* 0x0624 */;
            394: data_o = 32'h40878433 /* 0x0628 */;
            395: data_o = 32'h470186a2 /* 0x062c */;
            396: data_o = 32'hda7ff0ef /* 0x0630 */;
            397: data_o = 32'hb7e1d959 /* 0x0634 */;
            398: data_o = 32'h346dc7b7 /* 0x0638 */;
            399: data_o = 32'h5d678793 /* 0x063c */;
            400: data_o = 32'h38866737 /* 0x0640 */;
            401: data_o = 32'h94b70713 /* 0x0644 */;
            402: data_o = 32'h97ba1782 /* 0x0648 */;
            403: data_o = 32'h02f53833 /* 0x064c */;
            404: data_o = 32'h00040717 /* 0x0650 */;
            405: data_o = 32'h00040797 /* 0x0654 */;
            406: data_o = 32'h07136631 /* 0x0658 */;
            407: data_o = 32'h87939b07 /* 0x065c */;
            408: data_o = 32'h97329ac7 /* 0x0660 */;
            409: data_o = 32'h288397b2 /* 0x0664 */;
            410: data_o = 32'ha783ffc7 /* 0x0668 */;
            411: data_o = 32'h5813ff87 /* 0x066c */;
            412: data_o = 32'h18820098 /* 0x0670 */;
            413: data_o = 32'h93811782 /* 0x0674 */;
            414: data_o = 32'h00f8e8b3 /* 0x0678 */;
            415: data_o = 32'hb00025f3 /* 0x067c */;
            416: data_o = 32'h00040717 /* 0x0680 */;
            417: data_o = 32'h00040797 /* 0x0684 */;
            418: data_o = 32'h98070713 /* 0x0688 */;
            419: data_o = 32'h97c78793 /* 0x068c */;
            420: data_o = 32'h97b29732 /* 0x0690 */;
            421: data_o = 32'hffc72683 /* 0x0694 */;
            422: data_o = 32'hff87a783 /* 0x0698 */;
            423: data_o = 32'h17821682 /* 0x069c */;
            424: data_o = 32'h8edd9381 /* 0x06a0 */;
            425: data_o = 32'hfcd88ce3 /* 0x06a4 */;
            426: data_o = 32'h68b19836 /* 0x06a8 */;
            427: data_o = 32'hb0002373 /* 0x06ac */;
            428: data_o = 32'h00040717 /* 0x06b0 */;
            429: data_o = 32'h00040797 /* 0x06b4 */;
            430: data_o = 32'h95070713 /* 0x06b8 */;
            431: data_o = 32'h94c78793 /* 0x06bc */;
            432: data_o = 32'h974697c6 /* 0x06c0 */;
            433: data_o = 32'hffc72703 /* 0x06c4 */;
            434: data_o = 32'hff87a603 /* 0x06c8 */;
            435: data_o = 32'h02071793 /* 0x06cc */;
            436: data_o = 32'h02061713 /* 0x06d0 */;
            437: data_o = 32'h8fd99301 /* 0x06d4 */;
            438: data_o = 32'hfd07eae3 /* 0x06d8 */;
            439: data_o = 32'h40b30333 /* 0x06dc */;
            440: data_o = 32'h02a30533 /* 0x06e0 */;
            441: data_o = 32'h55338f95 /* 0x06e4 */;
            442: data_o = 32'h808202f5 /* 0x06e8 */;
            443: data_o = 32'h01002797 /* 0x06ec */;
            444: data_o = 32'h91478793 /* 0x06f0 */;
            445: data_o = 32'h0147c783 /* 0x06f4 */;
            446: data_o = 32'hcb898b85 /* 0x06f8 */;
            447: data_o = 32'h01002797 /* 0x06fc */;
            448: data_o = 32'h9047c503 /* 0x0700 */;
            449: data_o = 32'h35131569 /* 0x0704 */;
            450: data_o = 32'h80820015 /* 0x0708 */;
            451: data_o = 32'h80824501 /* 0x070c */;
            452: data_o = 32'h0733c585 /* 0x0710 */;
            453: data_o = 32'h279700b5 /* 0x0714 */;
            454: data_o = 32'h87930100 /* 0x0718 */;
            455: data_o = 32'hc7838ea7 /* 0x071c */;
            456: data_o = 32'h8b850147 /* 0x0720 */;
            457: data_o = 32'h2797dbed /* 0x0724 */;
            458: data_o = 32'hc7830100 /* 0x0728 */;
            459: data_o = 32'h05058da7 /* 0x072c */;
            460: data_o = 32'hfef50fa3 /* 0x0730 */;
            461: data_o = 32'hfee511e3 /* 0x0734 */;
            462: data_o = 32'h71798082 /* 0x0738 */;
            463: data_o = 32'hf022f406 /* 0x073c */;
            464: data_o = 32'h2797ec26 /* 0x0740 */;
            465: data_o = 32'h87930100 /* 0x0744 */;
            466: data_o = 32'hc7838be7 /* 0x0748 */;
            467: data_o = 32'hf7930147 /* 0x074c */;
            468: data_o = 32'hdbe50207 /* 0x0750 */;
            469: data_o = 32'h01002797 /* 0x0754 */;
            470: data_o = 32'h86234719 /* 0x0758 */;
            471: data_o = 32'h44c98ae7 /* 0x075c */;
            472: data_o = 32'h000f444d /* 0x0760 */;
            473: data_o = 32'h27970ff0 /* 0x0764 */;
            474: data_o = 32'h87930100 /* 0x0768 */;
            475: data_o = 32'hc78389a7 /* 0x076c */;
            476: data_o = 32'h8b850147 /* 0x0770 */;
            477: data_o = 32'h2797dbed /* 0x0774 */;
            478: data_o = 32'hc7830100 /* 0x0778 */;
            479: data_o = 32'hf71388a7 /* 0x077c */;
            480: data_o = 32'h85630ff7 /* 0x0780 */;
            481: data_o = 32'h00631097 /* 0x0784 */;
            482: data_o = 32'h47c50887 /* 0x0788 */;
            483: data_o = 32'h14f71963 /* 0x078c */;
            484: data_o = 32'h850a45a1 /* 0x0790 */;
            485: data_o = 32'hf7dff0ef /* 0x0794 */;
            486: data_o = 32'h45a10028 /* 0x0798 */;
            487: data_o = 32'hf75ff0ef /* 0x079c */;
            488: data_o = 32'h01002797 /* 0x07a0 */;
            489: data_o = 32'h86078793 /* 0x07a4 */;
            490: data_o = 32'h0147c783 /* 0x07a8 */;
            491: data_o = 32'h0207f793 /* 0x07ac */;
            492: data_o = 32'h6622dbe5 /* 0x07b0 */;
            493: data_o = 32'h27974719 /* 0x07b4 */;
            494: data_o = 32'h85230100 /* 0x07b8 */;
            495: data_o = 32'h670284e7 /* 0x07bc */;
            496: data_o = 32'h963ac605 /* 0x07c0 */;
            497: data_o = 32'h00074683 /* 0x07c4 */;
            498: data_o = 32'h01002797 /* 0x07c8 */;
            499: data_o = 32'h83878793 /* 0x07cc */;
            500: data_o = 32'h0147c783 /* 0x07d0 */;
            501: data_o = 32'h0207f793 /* 0x07d4 */;
            502: data_o = 32'h2797dbe5 /* 0x07d8 */;
            503: data_o = 32'h07050100 /* 0x07dc */;
            504: data_o = 32'h82d78323 /* 0x07e0 */;
            505: data_o = 32'hfec710e3 /* 0x07e4 */;
            506: data_o = 32'h01002797 /* 0x07e8 */;
            507: data_o = 32'h81878793 /* 0x07ec */;
            508: data_o = 32'h0147c783 /* 0x07f0 */;
            509: data_o = 32'h0207f793 /* 0x07f4 */;
            510: data_o = 32'h2797dbe5 /* 0x07f8 */;
            511: data_o = 32'h47110100 /* 0x07fc */;
            512: data_o = 32'h80e78323 /* 0x0800 */;
            513: data_o = 32'h45a1bfb9 /* 0x0804 */;
            514: data_o = 32'hf0ef850a /* 0x0808 */;
            515: data_o = 32'h1797f07f /* 0x080c */;
            516: data_o = 32'h87930100 /* 0x0810 */;
            517: data_o = 32'hc7837f27 /* 0x0814 */;
            518: data_o = 32'hf7930147 /* 0x0818 */;
            519: data_o = 32'hdbe50207 /* 0x081c */;
            520: data_o = 32'h01001797 /* 0x0820 */;
            521: data_o = 32'h80234719 /* 0x0824 */;
            522: data_o = 32'h000f7ee7 /* 0x0828 */;
            523: data_o = 32'h67820ff0 /* 0x082c */;
            524: data_o = 32'h0000100f /* 0x0830 */;
            525: data_o = 32'hc42a9782 /* 0x0834 */;
            526: data_o = 32'h0ff0000f /* 0x0838 */;
            527: data_o = 32'h01001797 /* 0x083c */;
            528: data_o = 32'h7c478793 /* 0x0840 */;
            529: data_o = 32'h0147c783 /* 0x0844 */;
            530: data_o = 32'h0207f793 /* 0x0848 */;
            531: data_o = 32'h4751dbe5 /* 0x084c */;
            532: data_o = 32'h01001797 /* 0x0850 */;
            533: data_o = 32'h7ae78823 /* 0x0854 */;
            534: data_o = 32'h00380070 /* 0x0858 */;
            535: data_o = 32'h00074683 /* 0x085c */;
            536: data_o = 32'h01001797 /* 0x0860 */;
            537: data_o = 32'h7a078793 /* 0x0864 */;
            538: data_o = 32'h0147c783 /* 0x0868 */;
            539: data_o = 32'h0207f793 /* 0x086c */;
            540: data_o = 32'h1797dbe5 /* 0x0870 */;
            541: data_o = 32'h07050100 /* 0x0874 */;
            542: data_o = 32'h78d78723 /* 0x0878 */;
            543: data_o = 32'hfee610e3 /* 0x087c */;
            544: data_o = 32'h70a24522 /* 0x0880 */;
            545: data_o = 32'h64e27402 /* 0x0884 */;
            546: data_o = 32'h80826145 /* 0x0888 */;
            547: data_o = 32'h850a45a1 /* 0x088c */;
            548: data_o = 32'he81ff0ef /* 0x0890 */;
            549: data_o = 32'h45a10028 /* 0x0894 */;
            550: data_o = 32'he79ff0ef /* 0x0898 */;
            551: data_o = 32'h01001797 /* 0x089c */;
            552: data_o = 32'h76478793 /* 0x08a0 */;
            553: data_o = 32'h0147c783 /* 0x08a4 */;
            554: data_o = 32'h0207f793 /* 0x08a8 */;
            555: data_o = 32'h65a2dbe5 /* 0x08ac */;
            556: data_o = 32'h17976502 /* 0x08b0 */;
            557: data_o = 32'h47190100 /* 0x08b4 */;
            558: data_o = 32'h74e78723 /* 0x08b8 */;
            559: data_o = 32'he55ff0ef /* 0x08bc */;
            560: data_o = 32'h01001797 /* 0x08c0 */;
            561: data_o = 32'h74078793 /* 0x08c4 */;
            562: data_o = 32'h0147c783 /* 0x08c8 */;
            563: data_o = 32'h0207f793 /* 0x08cc */;
            564: data_o = 32'h1797dbe5 /* 0x08d0 */;
            565: data_o = 32'h47110100 /* 0x08d4 */;
            566: data_o = 32'h72e78723 /* 0x08d8 */;
            567: data_o = 32'h4505b559 /* 0x08dc */;
            568: data_o = 32'hc93db74d /* 0x08e0 */;
            569: data_o = 32'h001c27b7 /* 0x08e4 */;
            570: data_o = 32'h02f55533 /* 0x08e8 */;
            571: data_o = 32'h01001717 /* 0x08ec */;
            572: data_o = 32'h71470713 /* 0x08f0 */;
            573: data_o = 32'h01001797 /* 0x08f4 */;
            574: data_o = 32'h00070223 /* 0x08f8 */;
            575: data_o = 32'h70c78793 /* 0x08fc */;
            576: data_o = 32'hf8000713 /* 0x0900 */;
            577: data_o = 32'h00e78623 /* 0x0904 */;
            578: data_o = 32'h01001597 /* 0x0908 */;
            579: data_o = 32'h01001617 /* 0x090c */;
            580: data_o = 32'h6f460613 /* 0x0910 */;
            581: data_o = 32'h01001697 /* 0x0914 */;
            582: data_o = 32'h6ec68693 /* 0x0918 */;
            583: data_o = 32'h1717430d /* 0x091c */;
            584: data_o = 32'h07130100 /* 0x0920 */;
            585: data_o = 32'h08936e27 /* 0x0924 */;
            586: data_o = 32'h1797fc70 /* 0x0928 */;
            587: data_o = 32'h87930100 /* 0x092c */;
            588: data_o = 32'h08136d67 /* 0x0930 */;
            589: data_o = 32'h7e130200 /* 0x0934 */;
            590: data_o = 32'h81210ff5 /* 0x0938 */;
            591: data_o = 32'h6fc58c23 /* 0x093c */;
            592: data_o = 32'h0ff57513 /* 0x0940 */;
            593: data_o = 32'h00a60223 /* 0x0944 */;
            594: data_o = 32'h00668623 /* 0x0948 */;
            595: data_o = 32'h01170423 /* 0x094c */;
            596: data_o = 32'h01078823 /* 0x0950 */;
            597: data_o = 32'h0ff0000f /* 0x0954 */;
            598: data_o = 32'h4e038082 /* 0x0958 */;
            599: data_o = 32'h43220001 /* 0x095c */;
            600: data_o = 32'hce31cd39 /* 0x0960 */;
            601: data_o = 32'h563bcda9 /* 0x0964 */;
            602: data_o = 32'h231902b6 /* 0x0968 */;
            603: data_o = 32'h131b65c1 /* 0x096c */;
            604: data_o = 32'h561b0023 /* 0x0970 */;
            605: data_o = 32'h367d0016 /* 0x0974 */;
            606: data_o = 32'h04b67363 /* 0x0978 */;
            607: data_o = 32'h01fe1e1b /* 0x097c */;
            608: data_o = 32'h01e8989b /* 0x0980 */;
            609: data_o = 32'h01c8e8b3 /* 0x0984 */;
            610: data_o = 32'h01d8181b /* 0x0988 */;
            611: data_o = 32'h68338bbd /* 0x098c */;
            612: data_o = 32'h979b0118 /* 0x0990 */;
            613: data_o = 32'h8b3d0187 /* 0x0994 */;
            614: data_o = 32'he7b3610c /* 0x0998 */;
            615: data_o = 32'h171b0107 /* 0x099c */;
            616: data_o = 32'h8abd0147 /* 0x09a0 */;
            617: data_o = 32'h13028f5d /* 0x09a4 */;
            618: data_o = 32'h0106969b /* 0x09a8 */;
            619: data_o = 32'h02035313 /* 0x09ac */;
            620: data_o = 32'h8ed18ed9 /* 0x09b0 */;
            621: data_o = 32'h006587b3 /* 0x09b4 */;
            622: data_o = 32'h4501c394 /* 0x09b8 */;
            623: data_o = 32'h450d8082 /* 0x09bc */;
            624: data_o = 32'h07b78082 /* 0x09c0 */;
            625: data_o = 32'hc91c4000 /* 0x09c4 */;
            626: data_o = 32'h9713495c /* 0x09c8 */;
            627: data_o = 32'h4de30217 /* 0x09cc */;
            628: data_o = 32'h4958fe07 /* 0x09d0 */;
            629: data_o = 32'h0087579b /* 0x09d4 */;
            630: data_o = 32'hf7938fd9 /* 0x09d8 */;
            631: data_o = 32'hfbf50ff7 /* 0x09dc */;
            632: data_o = 32'h00052823 /* 0x09e0 */;
            633: data_o = 32'hc9498082 /* 0x09e4 */;
            634: data_o = 32'he84a7179 /* 0x09e8 */;
            635: data_o = 32'h00853903 /* 0x09ec */;
            636: data_o = 32'hf406f022 /* 0x09f0 */;
            637: data_o = 32'h0f63842a /* 0x09f4 */;
            638: data_o = 32'hec260609 /* 0x09f8 */;
            639: data_o = 32'he26384ae /* 0x09fc */;
            640: data_o = 32'h35170725 /* 0x0a00 */;
            641: data_o = 32'h05130100 /* 0x0a04 */;
            642: data_o = 32'he0085fe5 /* 0x0a08 */;
            643: data_o = 32'hfb7ff0ef /* 0x0a0c */;
            644: data_o = 32'h470547bd /* 0x0a10 */;
            645: data_o = 32'h86bee43a /* 0x0a14 */;
            646: data_o = 32'he002873e /* 0x0a18 */;
            647: data_o = 32'h0004861b /* 0x0a1c */;
            648: data_o = 32'h0009059b /* 0x0a20 */;
            649: data_o = 32'h48818522 /* 0x0a24 */;
            650: data_o = 32'hf0ef4801 /* 0x0a28 */;
            651: data_o = 32'h87aaf31f /* 0x0a2c */;
            652: data_o = 32'hef9d450d /* 0x0a30 */;
            653: data_o = 32'h01003717 /* 0x0a34 */;
            654: data_o = 32'h5cc70713 /* 0x0a38 */;
            655: data_o = 32'h800006b7 /* 0x0a3c */;
            656: data_o = 32'h01003797 /* 0x0a40 */;
            657: data_o = 32'h8793cb14 /* 0x0a44 */;
            658: data_o = 32'h4b985c07 /* 0x0a48 */;
            659: data_o = 32'h200006b7 /* 0x0a4c */;
            660: data_o = 32'h01003797 /* 0x0a50 */;
            661: data_o = 32'h87938f55 /* 0x0a54 */;
            662: data_o = 32'h64e25b07 /* 0x0a58 */;
            663: data_o = 32'h4501cb98 /* 0x0a5c */;
            664: data_o = 32'h64e2a019 /* 0x0a60 */;
            665: data_o = 32'h70a24551 /* 0x0a64 */;
            666: data_o = 32'h69427402 /* 0x0a68 */;
            667: data_o = 32'h80826145 /* 0x0a6c */;
            668: data_o = 32'hbfd564e2 /* 0x0a70 */;
            669: data_o = 32'hbfc5454d /* 0x0a74 */;
            670: data_o = 32'h80824545 /* 0x0a78 */;
            671: data_o = 32'he0221141 /* 0x0a7c */;
            672: data_o = 32'h0437e406 /* 0x0a80 */;
            673: data_o = 32'hf0ef0300 /* 0x0a84 */;
            674: data_o = 32'h0793e5df /* 0x0a88 */;
            675: data_o = 32'h47980004 /* 0x0a8c */;
            676: data_o = 32'hcf198b09 /* 0x0a90 */;
            677: data_o = 32'h0007a423 /* 0x0a94 */;
            678: data_o = 32'h278343c8 /* 0x0a98 */;
            679: data_o = 32'h64020004 /* 0x0a9c */;
            680: data_o = 32'h178260a2 /* 0x0aa0 */;
            681: data_o = 32'h93811502 /* 0x0aa4 */;
            682: data_o = 32'h01418d5d /* 0x0aa8 */;
            683: data_o = 32'he0cff06f /* 0x0aac */;
            684: data_o = 32'hc3dff0ef /* 0x0ab0 */;
            685: data_o = 32'h6402d979 /* 0x0ab4 */;
            686: data_o = 32'h014160a2 /* 0x0ab8 */;
            687: data_o = 32'h7119b9bd /* 0x0abc */;
            688: data_o = 32'hf4a6f8a2 /* 0x0ac0 */;
            689: data_o = 32'hf0cafc86 /* 0x0ac4 */;
            690: data_o = 32'h842eecce /* 0x0ac8 */;
            691: data_o = 32'h46a184aa /* 0x0acc */;
            692: data_o = 32'h0613852e /* 0x0ad0 */;
            693: data_o = 32'h100c2000 /* 0x0ad4 */;
            694: data_o = 32'hed799482 /* 0x0ad8 */;
            695: data_o = 32'h545247b7 /* 0x0adc */;
            696: data_o = 32'h15078793 /* 0x0ae0 */;
            697: data_o = 32'h20494737 /* 0x0ae4 */;
            698: data_o = 32'h17827682 /* 0x0ae8 */;
            699: data_o = 32'h64570713 /* 0x0aec */;
            700: data_o = 32'h936397ba /* 0x0af0 */;
            701: data_o = 32'h46c10cf6 /* 0x0af4 */;
            702: data_o = 32'h24800613 /* 0x0af8 */;
            703: data_o = 32'h8522858a /* 0x0afc */;
            704: data_o = 32'h87aa9482 /* 0x0b00 */;
            705: data_o = 32'h12051563 /* 0x0b04 */;
            706: data_o = 32'hc7dd47a2 /* 0x0b08 */;
            707: data_o = 32'he0dae4d6 /* 0x0b0c */;
            708: data_o = 32'h4ce50ab7 /* 0x0b10 */;
            709: data_o = 32'h622c4b37 /* 0x0b14 */;
            710: data_o = 32'hd95a8a93 /* 0x0b18 */;
            711: data_o = 32'h0269b737 /* 0x0b1c */;
            712: data_o = 32'h101b0b13 /* 0x0b20 */;
            713: data_o = 32'h1494d7b7 /* 0x0b24 */;
            714: data_o = 32'h07131a82 /* 0x0b28 */;
            715: data_o = 32'h1b0226a7 /* 0x0b2c */;
            716: data_o = 32'hf9878793 /* 0x0b30 */;
            717: data_o = 32'h05f00913 /* 0x0b34 */;
            718: data_o = 32'hf862e8d2 /* 0x0b38 */;
            719: data_o = 32'h9abafc5e /* 0x0b3c */;
            720: data_o = 32'h8a4a9b3e /* 0x0b40 */;
            721: data_o = 32'h4c014981 /* 0x0b44 */;
            722: data_o = 32'h00c16783 /* 0x0b48 */;
            723: data_o = 32'h46c16b82 /* 0x0b4c */;
            724: data_o = 32'h038787b3 /* 0x0b50 */;
            725: data_o = 32'h05b30ba6 /* 0x0b54 */;
            726: data_o = 32'h852200d1 /* 0x0b58 */;
            727: data_o = 32'h86139bbe /* 0x0b5c */;
            728: data_o = 32'h9482020b /* 0x0b60 */;
            729: data_o = 32'h46c187aa /* 0x0b64 */;
            730: data_o = 32'h100c865e /* 0x0b68 */;
            731: data_o = 32'hebdd8522 /* 0x0b6c */;
            732: data_o = 32'h67e26742 /* 0x0b70 */;
            733: data_o = 32'h000c1863 /* 0x0b74 */;
            734: data_o = 32'h05f70913 /* 0x0b78 */;
            735: data_o = 32'h0127f363 /* 0x0b7c */;
            736: data_o = 32'h89ba893e /* 0x0b80 */;
            737: data_o = 32'h68638f99 /* 0x0b84 */;
            738: data_o = 32'h948200fa /* 0x0b88 */;
            739: data_o = 32'he95987aa /* 0x0b8c */;
            740: data_o = 32'h85637782 /* 0x0b90 */;
            741: data_o = 32'h67830957 /* 0x0b94 */;
            742: data_o = 32'h0c050081 /* 0x0b98 */;
            743: data_o = 32'hfafc46e3 /* 0x0b9c */;
            744: data_o = 32'h00816783 /* 0x0ba0 */;
            745: data_o = 32'h01878463 /* 0x0ba4 */;
            746: data_o = 32'h696269c2 /* 0x0ba8 */;
            747: data_o = 32'h6aa66a46 /* 0x0bac */;
            748: data_o = 32'h7be26b06 /* 0x0bb0 */;
            749: data_o = 32'ha0217c42 /* 0x0bb4 */;
            750: data_o = 32'h05f00913 /* 0x0bb8 */;
            751: data_o = 32'h06934981 /* 0x0bbc */;
            752: data_o = 32'h86b30019 /* 0x0bc0 */;
            753: data_o = 32'hf5974136 /* 0x0bc4 */;
            754: data_o = 32'h06a60dff /* 0x0bc8 */;
            755: data_o = 32'h00999613 /* 0x0bcc */;
            756: data_o = 32'h43a58593 /* 0x0bd0 */;
            757: data_o = 32'h94828522 /* 0x0bd4 */;
            758: data_o = 32'he93187aa /* 0x0bd8 */;
            759: data_o = 32'h0014e493 /* 0x0bdc */;
            760: data_o = 32'hf7172481 /* 0x0be0 */;
            761: data_o = 32'hf79700ff /* 0x0be4 */;
            762: data_o = 32'h240100ff /* 0x0be8 */;
            763: data_o = 32'h40972f23 /* 0x0bec */;
            764: data_o = 32'h41a78793 /* 0x0bf0 */;
            765: data_o = 32'h870ec3c0 /* 0x0bf4 */;
            766: data_o = 32'h00fff797 /* 0x0bf8 */;
            767: data_o = 32'h70e67446 /* 0x0bfc */;
            768: data_o = 32'h790674a6 /* 0x0c00 */;
            769: data_o = 32'h270169e6 /* 0x0c04 */;
            770: data_o = 32'h40878793 /* 0x0c08 */;
            771: data_o = 32'h0dfff517 /* 0x0c0c */;
            772: data_o = 32'h0513c7d8 /* 0x0c10 */;
            773: data_o = 32'h61093f45 /* 0x0c14 */;
            774: data_o = 32'hca0ff06f /* 0x0c18 */;
            775: data_o = 32'h9ce377a2 /* 0x0c1c */;
            776: data_o = 32'hbfbdf767 /* 0x0c20 */;
            777: data_o = 32'h6aa66a46 /* 0x0c24 */;
            778: data_o = 32'h7be26b06 /* 0x0c28 */;
            779: data_o = 32'h70e67c42 /* 0x0c2c */;
            780: data_o = 32'h74a67446 /* 0x0c30 */;
            781: data_o = 32'h69e67906 /* 0x0c34 */;
            782: data_o = 32'h6109853e /* 0x0c38 */;
            783: data_o = 32'h09638082 /* 0x0c3c */;
            784: data_o = 32'h87631605 /* 0x0c40 */;
            785: data_o = 32'h11411605 /* 0x0c44 */;
            786: data_o = 32'he402e002 /* 0x0c48 */;
            787: data_o = 32'h0035f793 /* 0x0c4c */;
            788: data_o = 32'h6841cb9d /* 0x0c50 */;
            789: data_o = 32'hf0080813 /* 0x0c54 */;
            790: data_o = 32'h03138e0a /* 0x0c58 */;
            791: data_o = 32'hca590041 /* 0x0c5c */;
            792: data_o = 32'h5d634702 /* 0x0c60 */;
            793: data_o = 32'h377d0ae0 /* 0x0c64 */;
            794: data_o = 32'h00814683 /* 0x0c68 */;
            795: data_o = 32'h367d67a2 /* 0x0c6c */;
            796: data_o = 32'h00d58023 /* 0x0c70 */;
            797: data_o = 32'h058583a1 /* 0x0c74 */;
            798: data_o = 32'h1642e43e /* 0x0c78 */;
            799: data_o = 32'hf793c03a /* 0x0c7c */;
            800: data_o = 32'h92410035 /* 0x0c80 */;
            801: data_o = 32'h430dffe9 /* 0x0c84 */;
            802: data_o = 32'h7e6386ae /* 0x0c88 */;
            803: data_o = 32'h66c102c3 /* 0x0c8c */;
            804: data_o = 32'h079b16f1 /* 0x0c90 */;
            805: data_o = 32'h4702ffc6 /* 0x0c94 */;
            806: data_o = 32'h68c18ff5 /* 0x0c98 */;
            807: data_o = 32'h00458693 /* 0x0c9c */;
            808: data_o = 32'h889396be /* 0x0ca0 */;
            809: data_o = 32'h8f0af008 /* 0x0ca4 */;
            810: data_o = 32'h00410e93 /* 0x0ca8 */;
            811: data_o = 32'h04e35663 /* 0x0cac */;
            812: data_o = 32'h48223771 /* 0x0cb0 */;
            813: data_o = 32'hc03a47b2 /* 0x0cb4 */;
            814: data_o = 32'h0105a023 /* 0x0cb8 */;
            815: data_o = 32'h0591c43e /* 0x0cbc */;
            816: data_o = 32'hfeb696e3 /* 0x0cc0 */;
            817: data_o = 32'hc61d8a0d /* 0x0cc4 */;
            818: data_o = 32'h87b69e35 /* 0x0cc8 */;
            819: data_o = 32'h16424682 /* 0x0ccc */;
            820: data_o = 32'h5d639241 /* 0x0cd0 */;
            821: data_o = 32'h36fd08d0 /* 0x0cd4 */;
            822: data_o = 32'h00814583 /* 0x0cd8 */;
            823: data_o = 32'h07856722 /* 0x0cdc */;
            824: data_o = 32'hfeb78fa3 /* 0x0ce0 */;
            825: data_o = 32'h95938321 /* 0x0ce4 */;
            826: data_o = 32'hc0360307 /* 0x0ce8 */;
            827: data_o = 32'he43a91c1 /* 0x0cec */;
            828: data_o = 32'hfec591e3 /* 0x0cf0 */;
            829: data_o = 32'h80820141 /* 0x0cf4 */;
            830: data_o = 32'h00053803 /* 0x0cf8 */;
            831: data_o = 32'h01482783 /* 0x0cfc */;
            832: data_o = 32'h0117f7b3 /* 0x0d00 */;
            833: data_o = 32'h2783dfe5 /* 0x0d04 */;
            834: data_o = 32'h781302c8 /* 0x0d08 */;
            835: data_o = 32'h27810037 /* 0x0d0c */;
            836: data_o = 32'h02081563 /* 0x0d10 */;
            837: data_o = 32'hc71c970a /* 0x0d14 */;
            838: data_o = 32'hbf614702 /* 0x0d18 */;
            839: data_o = 32'h4adc6114 /* 0x0d1c */;
            840: data_o = 32'h0107f7b3 /* 0x0d20 */;
            841: data_o = 32'h56dcdfed /* 0x0d24 */;
            842: data_o = 32'h00377693 /* 0x0d28 */;
            843: data_o = 32'he2952781 /* 0x0d2c */;
            844: data_o = 32'hc71c970a /* 0x0d30 */;
            845: data_o = 32'h270d4702 /* 0x0d34 */;
            846: data_o = 32'h0833bf05 /* 0x0d38 */;
            847: data_o = 32'h8e3301e7 /* 0x0d3c */;
            848: data_o = 32'h042300ee /* 0x0d40 */;
            849: data_o = 32'h080500f8 /* 0x0d44 */;
            850: data_o = 32'h0087d79b /* 0x0d48 */;
            851: data_o = 32'hffc81be3 /* 0x0d4c */;
            852: data_o = 32'h06b3b78d /* 0x0d50 */;
            853: data_o = 32'h08b301c7 /* 0x0d54 */;
            854: data_o = 32'h842300e3 /* 0x0d58 */;
            855: data_o = 32'h068500f6 /* 0x0d5c */;
            856: data_o = 32'h0087d79b /* 0x0d60 */;
            857: data_o = 32'hff169be3 /* 0x0d64 */;
            858: data_o = 32'hbdfd270d /* 0x0d68 */;
            859: data_o = 32'h00053803 /* 0x0d6c */;
            860: data_o = 32'h859365c1 /* 0x0d70 */;
            861: data_o = 32'h2703f005 /* 0x0d74 */;
            862: data_o = 32'h8f6d0148 /* 0x0d78 */;
            863: data_o = 32'h2583df6d /* 0x0d7c */;
            864: data_o = 32'hf71302c8 /* 0x0d80 */;
            865: data_o = 32'h25810036 /* 0x0d84 */;
            866: data_o = 32'h0813cf19 /* 0x0d88 */;
            867: data_o = 32'h07330041 /* 0x0d8c */;
            868: data_o = 32'h983600d1 /* 0x0d90 */;
            869: data_o = 32'h00b70423 /* 0x0d94 */;
            870: data_o = 32'hd59b0705 /* 0x0d98 */;
            871: data_o = 32'h1be30085 /* 0x0d9c */;
            872: data_o = 32'h268dff07 /* 0x0da0 */;
            873: data_o = 32'h968abf15 /* 0x0da4 */;
            874: data_o = 32'h4682c68c /* 0x0da8 */;
            875: data_o = 32'hb72d268d /* 0x0dac */;
            876: data_o = 32'hcd418082 /* 0x0db0 */;
            877: data_o = 32'hf793c9d9 /* 0x0db4 */;
            878: data_o = 32'h06930035 /* 0x0db8 */;
            879: data_o = 32'hc39d0480 /* 0x0dbc */;
            880: data_o = 32'h6118c651 /* 0x0dc0 */;
            881: data_o = 32'hf7934b5c /* 0x0dc4 */;
            882: data_o = 32'h8de30ff7 /* 0x0dc8 */;
            883: data_o = 32'hc783fed7 /* 0x0dcc */;
            884: data_o = 32'h367d0005 /* 0x0dd0 */;
            885: data_o = 32'h08230585 /* 0x0dd4 */;
            886: data_o = 32'h164202f7 /* 0x0dd8 */;
            887: data_o = 32'h0035f793 /* 0x0ddc */;
            888: data_o = 32'hfff99241 /* 0x0de0 */;
            889: data_o = 32'h882e478d /* 0x0de4 */;
            890: data_o = 32'h02c7f963 /* 0x0de8 */;
            891: data_o = 32'h17f167c1 /* 0x0dec */;
            892: data_o = 32'hffc6081b /* 0x0df0 */;
            893: data_o = 32'h78336118 /* 0x0df4 */;
            894: data_o = 32'h879300f8 /* 0x0df8 */;
            895: data_o = 32'h983e0045 /* 0x0dfc */;
            896: data_o = 32'h04800693 /* 0x0e00 */;
            897: data_o = 32'hf7934b5c /* 0x0e04 */;
            898: data_o = 32'h8de30ff7 /* 0x0e08 */;
            899: data_o = 32'h419cfed7 /* 0x0e0c */;
            900: data_o = 32'hdb1c0591 /* 0x0e10 */;
            901: data_o = 32'hff0598e3 /* 0x0e14 */;
            902: data_o = 32'hca058a0d /* 0x0e18 */;
            903: data_o = 32'h00c8073b /* 0x0e1c */;
            904: data_o = 32'h85c21742 /* 0x0e20 */;
            905: data_o = 32'h06139341 /* 0x0e24 */;
            906: data_o = 32'h61140480 /* 0x0e28 */;
            907: data_o = 32'hf7934adc /* 0x0e2c */;
            908: data_o = 32'h8de30ff7 /* 0x0e30 */;
            909: data_o = 32'hc803fec7 /* 0x0e34 */;
            910: data_o = 32'h05850005 /* 0x0e38 */;
            911: data_o = 32'h03059793 /* 0x0e3c */;
            912: data_o = 32'h882393c1 /* 0x0e40 */;
            913: data_o = 32'h92e30306 /* 0x0e44 */;
            914: data_o = 32'h8082fee7 /* 0x0e48 */;
            915: data_o = 32'h41948082 /* 0x0e4c */;
            916: data_o = 32'hf0227179 /* 0x0e50 */;
            917: data_o = 32'hf406e44e /* 0x0e54 */;
            918: data_o = 32'he84aec26 /* 0x0e58 */;
            919: data_o = 32'h87ae4711 /* 0x0e5c */;
            920: data_o = 32'h89aa8432 /* 0x0e60 */;
            921: data_o = 32'h06e68863 /* 0x0e64 */;
            922: data_o = 32'h8b634715 /* 0x0e68 */;
            923: data_o = 32'h470d04e6 /* 0x0e6c */;
            924: data_o = 32'h06e69863 /* 0x0e70 */;
            925: data_o = 32'h0185d483 /* 0x0e74 */;
            926: data_o = 32'ha903698c /* 0x0e78 */;
            927: data_o = 32'h86260087 /* 0x0e7c */;
            928: data_o = 32'hf33ff0ef /* 0x0e80 */;
            929: data_o = 32'h44136709 /* 0x0e84 */;
            930: data_o = 32'h67850014 /* 0x0e88 */;
            931: data_o = 32'h0094141b /* 0x0e8c */;
            932: data_o = 32'h00a9191b /* 0x0e90 */;
            933: data_o = 32'hc0078793 /* 0x0e94 */;
            934: data_o = 32'h79338c59 /* 0x0e98 */;
            935: data_o = 32'hb70300f9 /* 0x0e9c */;
            936: data_o = 32'h34fd0009 /* 0x0ea0 */;
            937: data_o = 32'h1ff4f493 /* 0x0ea4 */;
            938: data_o = 32'h01246433 /* 0x0ea8 */;
            939: data_o = 32'h70a28c45 /* 0x0eac */;
            940: data_o = 32'h7402d700 /* 0x0eb0 */;
            941: data_o = 32'h694264e2 /* 0x0eb4 */;
            942: data_o = 32'h450169a2 /* 0x0eb8 */;
            943: data_o = 32'h80826145 /* 0x0ebc */;
            944: data_o = 32'h0205d483 /* 0x0ec0 */;
            945: data_o = 32'ha903698c /* 0x0ec4 */;
            946: data_o = 32'h86260087 /* 0x0ec8 */;
            947: data_o = 32'hee7ff0ef /* 0x0ecc */;
            948: data_o = 32'hbf55670d /* 0x0ed0 */;
            949: data_o = 32'h0085a903 /* 0x0ed4 */;
            950: data_o = 32'h0185d483 /* 0x0ed8 */;
            951: data_o = 32'hb7656705 /* 0x0edc */;
            952: data_o = 32'h740270a2 /* 0x0ee0 */;
            953: data_o = 32'h694264e2 /* 0x0ee4 */;
            954: data_o = 32'h853a69a2 /* 0x0ee8 */;
            955: data_o = 32'h80826145 /* 0x0eec */;
            956: data_o = 32'he8221101 /* 0x0ef0 */;
            957: data_o = 32'he04ae426 /* 0x0ef4 */;
            958: data_o = 32'h842aec06 /* 0x0ef8 */;
            959: data_o = 32'h84b2892e /* 0x0efc */;
            960: data_o = 32'h04800713 /* 0x0f00 */;
            961: data_o = 32'hf793485c /* 0x0f04 */;
            962: data_o = 32'h8de30ff7 /* 0x0f08 */;
            963: data_o = 32'h2503fee7 /* 0x0f0c */;
            964: data_o = 32'hf0ef0109 /* 0x0f10 */;
            965: data_o = 32'h2703a6cf /* 0x0f14 */;
            966: data_o = 32'h478500c9 /* 0x0f18 */;
            967: data_o = 32'h02f70d63 /* 0x0f1c */;
            968: data_o = 32'h0085551b /* 0x0f20 */;
            969: data_o = 32'h4689d808 /* 0x0f24 */;
            970: data_o = 32'h00892783 /* 0x0f28 */;
            971: data_o = 32'h0014c493 /* 0x0f2c */;
            972: data_o = 32'h07136705 /* 0x0f30 */;
            973: data_o = 32'h979bc007 /* 0x0f34 */;
            974: data_o = 32'h949b00a7 /* 0x0f38 */;
            975: data_o = 32'h8cd50094 /* 0x0f3c */;
            976: data_o = 32'h8fc58ff9 /* 0x0f40 */;
            977: data_o = 32'h8fd96709 /* 0x0f44 */;
            978: data_o = 32'hd41c60e2 /* 0x0f48 */;
            979: data_o = 32'h64a26442 /* 0x0f4c */;
            980: data_o = 32'h61056902 /* 0x0f50 */;
            981: data_o = 32'hd8088082 /* 0x0f54 */;
            982: data_o = 32'hb7f9468d /* 0x0f58 */;
            983: data_o = 32'h6118495c /* 0x0f5c */;
            984: data_o = 32'h4b5cd35c /* 0x0f60 */;
            985: data_o = 32'h01f7d79b /* 0x0f64 */;
            986: data_o = 32'h479ddfed /* 0x0f68 */;
            987: data_o = 32'h4501d71c /* 0x0f6c */;
            988: data_o = 32'h71518082 /* 0x0f70 */;
            989: data_o = 32'h8b2af95a /* 0x0f74 */;
            990: data_o = 32'hf7b76508 /* 0x0f78 */;
            991: data_o = 32'hf58602fa /* 0x0f7c */;
            992: data_o = 32'h07f78793 /* 0x0f80 */;
            993: data_o = 32'h1aa7e563 /* 0x0f84 */;
            994: data_o = 32'hf55eeda6 /* 0x0f88 */;
            995: data_o = 32'h4b8184b6 /* 0x0f8c */;
            996: data_o = 32'h10068163 /* 0x0f90 */;
            997: data_o = 32'he9caf1a2 /* 0x0f94 */;
            998: data_o = 32'he1d2e5ce /* 0x0f98 */;
            999: data_o = 32'hf162fd56 /* 0x0f9c */;
            1000: data_o = 32'he96aed66 /* 0x0fa0 */;
            1001: data_o = 32'h8a2ee56e /* 0x0fa4 */;
            1002: data_o = 32'h49858ab2 /* 0x0fa8 */;
            1003: data_o = 32'h440d4911 /* 0x0fac */;
            1004: data_o = 32'h017a87bb /* 0x0fb0 */;
            1005: data_o = 32'h017a0633 /* 0x0fb4 */;
            1006: data_o = 32'hf802e802 /* 0x0fb8 */;
            1007: data_o = 32'he082fc02 /* 0x0fbc */;
            1008: data_o = 32'h474dec82 /* 0x0fc0 */;
            1009: data_o = 32'hf4b2c0be /* 0x0fc4 */;
            1010: data_o = 32'hec02e402 /* 0x0fc8 */;
            1011: data_o = 32'hf402f002 /* 0x0fcc */;
            1012: data_o = 32'he882e482 /* 0x0fd0 */;
            1013: data_o = 32'hfc82f082 /* 0x0fd4 */;
            1014: data_o = 32'h00e10823 /* 0x0fd8 */;
            1015: data_o = 32'hde4ed84e /* 0x0fdc */;
            1016: data_o = 32'h87b3ccca /* 0x0fe0 */;
            1017: data_o = 32'h06134174 /* 0x0fe4 */;
            1018: data_o = 32'h73631000 /* 0x0fe8 */;
            1019: data_o = 32'h87b200f6 /* 0x0fec */;
            1020: data_o = 32'h010b2603 /* 0x0ff0 */;
            1021: data_o = 32'h000b3503 /* 0x0ff4 */;
            1022: data_o = 32'h00810d93 /* 0x0ff8 */;
            1023: data_o = 32'hd150f8be /* 0x0ffc */;
            1024: data_o = 32'h4c018cee /* 0x1000 */;
            1025: data_o = 32'h06134d09 /* 0x1004 */;
            1026: data_o = 32'h3613ffec /* 0x1008 */;
            1027: data_o = 32'h495c0016 /* 0x100c */;
            1028: data_o = 32'h01f7d79b /* 0x1010 */;
            1029: data_o = 32'ha783dfed /* 0x1014 */;
            1030: data_o = 32'h8263000c /* 0x1018 */;
            1031: data_o = 32'h61630fa7 /* 0x101c */;
            1032: data_o = 32'hc7dd08fd /* 0x1020 */;
            1033: data_o = 32'hf0ef85e6 /* 0x1024 */;
            1034: data_o = 32'h0c05ecbf /* 0x1028 */;
            1035: data_o = 32'h028c8c93 /* 0x102c */;
            1036: data_o = 32'h028c0463 /* 0x1030 */;
            1037: data_o = 32'h000b3503 /* 0x1034 */;
            1038: data_o = 32'h4715b7f9 /* 0x1038 */;
            1039: data_o = 32'h9863855a /* 0x103c */;
            1040: data_o = 32'hd60300e7 /* 0x1040 */;
            1041: data_o = 32'hb583020d /* 0x1044 */;
            1042: data_o = 32'hf0ef018d /* 0x1048 */;
            1043: data_o = 32'h8d93bf5f /* 0x104c */;
            1044: data_o = 32'h011c028d /* 0x1050 */;
            1045: data_o = 32'h03b78263 /* 0x1054 */;
            1046: data_o = 32'h000da783 /* 0x1058 */;
            1047: data_o = 32'hfd279fe3 /* 0x105c */;
            1048: data_o = 32'h018dd603 /* 0x1060 */;
            1049: data_o = 32'h010db583 /* 0x1064 */;
            1050: data_o = 32'h8d93855a /* 0x1068 */;
            1051: data_o = 32'hf0ef028d /* 0x106c */;
            1052: data_o = 32'h011cbd1f /* 0x1070 */;
            1053: data_o = 32'hffb792e3 /* 0x1074 */;
            1054: data_o = 32'h100b8b93 /* 0x1078 */;
            1055: data_o = 32'hf29beae3 /* 0x107c */;
            1056: data_o = 32'h694e740e /* 0x1080 */;
            1057: data_o = 32'h6a0e69ae /* 0x1084 */;
            1058: data_o = 32'h7c0a7aea /* 0x1088 */;
            1059: data_o = 32'h6d4a6cea /* 0x108c */;
            1060: data_o = 32'h70ae6daa /* 0x1090 */;
            1061: data_o = 32'h7baa64ee /* 0x1094 */;
            1062: data_o = 32'h45017b4a /* 0x1098 */;
            1063: data_o = 32'h8082616d /* 0x109c */;
            1064: data_o = 32'h676337f5 /* 0x10a0 */;
            1065: data_o = 32'h85e600fd /* 0x10a4 */;
            1066: data_o = 32'hf0ef855a /* 0x10a8 */;
            1067: data_o = 32'hdd35da5f /* 0x10ac */;
            1068: data_o = 32'h70ae740e /* 0x10b0 */;
            1069: data_o = 32'h694e64ee /* 0x10b4 */;
            1070: data_o = 32'h6a0e69ae /* 0x10b8 */;
            1071: data_o = 32'h7baa7aea /* 0x10bc */;
            1072: data_o = 32'h6cea7c0a /* 0x10c0 */;
            1073: data_o = 32'h6daa6d4a /* 0x10c4 */;
            1074: data_o = 32'h450d7b4a /* 0x10c8 */;
            1075: data_o = 32'h8082616d /* 0x10cc */;
            1076: data_o = 32'h04800613 /* 0x10d0 */;
            1077: data_o = 32'hf793495c /* 0x10d4 */;
            1078: data_o = 32'h8de30ff7 /* 0x10d8 */;
            1079: data_o = 32'hc603fec7 /* 0x10dc */;
            1080: data_o = 32'h0793008c /* 0x10e0 */;
            1081: data_o = 32'h37b3ffec /* 0x10e4 */;
            1082: data_o = 32'h082300f0 /* 0x10e8 */;
            1083: data_o = 32'h360302c5 /* 0x10ec */;
            1084: data_o = 32'h979b000b /* 0x10f0 */;
            1085: data_o = 32'h65890097 /* 0x10f4 */;
            1086: data_o = 32'hd61c8fcd /* 0x10f8 */;
            1087: data_o = 32'ha583b73d /* 0x10fc */;
            1088: data_o = 32'hd603008c /* 0x1100 */;
            1089: data_o = 32'h6805010c /* 0x1104 */;
            1090: data_o = 32'hffec0793 /* 0x1108 */;
            1091: data_o = 32'h00a5959b /* 0x110c */;
            1092: data_o = 32'hc0080813 /* 0x1110 */;
            1093: data_o = 32'h00f037b3 /* 0x1114 */;
            1094: data_o = 32'h0105f5b3 /* 0x1118 */;
            1095: data_o = 32'h0097979b /* 0x111c */;
            1096: data_o = 32'h8fcd367d /* 0x1120 */;
            1097: data_o = 32'h1ff67613 /* 0x1124 */;
            1098: data_o = 32'hd51c8fd1 /* 0x1128 */;
            1099: data_o = 32'h70aebdfd /* 0x112c */;
            1100: data_o = 32'h45557b4a /* 0x1130 */;
            1101: data_o = 32'h8082616d /* 0x1134 */;
            1102: data_o = 32'he4261101 /* 0x1138 */;
            1103: data_o = 32'h610884aa /* 0x113c */;
            1104: data_o = 32'hec06e822 /* 0x1140 */;
            1105: data_o = 32'hd14c8432 /* 0x1144 */;
            1106: data_o = 32'hd79b495c /* 0x1148 */;
            1107: data_o = 32'hdfed01f7 /* 0x114c */;
            1108: data_o = 32'h4709401c /* 0x1150 */;
            1109: data_o = 32'h06e78663 /* 0x1154 */;
            1110: data_o = 32'h02f76463 /* 0x1158 */;
            1111: data_o = 32'h4601c3a9 /* 0x115c */;
            1112: data_o = 32'hf0ef85a2 /* 0x1160 */;
            1113: data_o = 32'h4018d8ff /* 0x1164 */;
            1114: data_o = 32'h04634791 /* 0x1168 */;
            1115: data_o = 32'h479508f7 /* 0x116c */;
            1116: data_o = 32'h06f70963 /* 0x1170 */;
            1117: data_o = 32'h60e24501 /* 0x1174 */;
            1118: data_o = 32'h64a26442 /* 0x1178 */;
            1119: data_o = 32'h80826105 /* 0x117c */;
            1120: data_o = 32'h686337f5 /* 0x1180 */;
            1121: data_o = 32'h460100f7 /* 0x1184 */;
            1122: data_o = 32'h852685a2 /* 0x1188 */;
            1123: data_o = 32'hcc3ff0ef /* 0x118c */;
            1124: data_o = 32'h60e2d979 /* 0x1190 */;
            1125: data_o = 32'h64a26442 /* 0x1194 */;
            1126: data_o = 32'h6105450d /* 0x1198 */;
            1127: data_o = 32'h07138082 /* 0x119c */;
            1128: data_o = 32'h495c0480 /* 0x11a0 */;
            1129: data_o = 32'h0ff7f793 /* 0x11a4 */;
            1130: data_o = 32'hfee78de3 /* 0x11a8 */;
            1131: data_o = 32'h00844703 /* 0x11ac */;
            1132: data_o = 32'h87936789 /* 0x11b0 */;
            1133: data_o = 32'h08232007 /* 0x11b4 */;
            1134: data_o = 32'h609802e5 /* 0x11b8 */;
            1135: data_o = 32'hb765d71c /* 0x11bc */;
            1136: data_o = 32'h01045783 /* 0x11c0 */;
            1137: data_o = 32'h66854418 /* 0x11c4 */;
            1138: data_o = 32'h171b37fd /* 0x11c8 */;
            1139: data_o = 32'h869300a7 /* 0x11cc */;
            1140: data_o = 32'hf793c006 /* 0x11d0 */;
            1141: data_o = 32'h8f751ff7 /* 0x11d4 */;
            1142: data_o = 32'he7938fd9 /* 0x11d8 */;
            1143: data_o = 32'hd51c2007 /* 0x11dc */;
            1144: data_o = 32'h5603b759 /* 0x11e0 */;
            1145: data_o = 32'h6c0c0204 /* 0x11e4 */;
            1146: data_o = 32'hf0ef8526 /* 0x11e8 */;
            1147: data_o = 32'h4501a55f /* 0x11ec */;
            1148: data_o = 32'h5603b759 /* 0x11f0 */;
            1149: data_o = 32'h680c0184 /* 0x11f4 */;
            1150: data_o = 32'hf0ef8526 /* 0x11f8 */;
            1151: data_o = 32'h4501a45f /* 0x11fc */;
            1152: data_o = 32'h7119bf9d /* 0x1200 */;
            1153: data_o = 32'hf0caf8a2 /* 0x1204 */;
            1154: data_o = 32'he0dae4d6 /* 0x1208 */;
            1155: data_o = 32'he42efc86 /* 0x120c */;
            1156: data_o = 32'h8b32842a /* 0x1210 */;
            1157: data_o = 32'h8aba8936 /* 0x1214 */;
            1158: data_o = 32'h0793cdb1 /* 0x1218 */;
            1159: data_o = 32'h80630fd0 /* 0x121c */;
            1160: data_o = 32'h469912f5 /* 0x1220 */;
            1161: data_o = 32'h470d480c /* 0x1224 */;
            1162: data_o = 32'h0830003c /* 0x1228 */;
            1163: data_o = 32'hce028522 /* 0x122c */;
            1164: data_o = 32'hd202d002 /* 0x1230 */;
            1165: data_o = 32'hde02dc02 /* 0x1234 */;
            1166: data_o = 32'hcc3af836 /* 0x1238 */;
            1167: data_o = 32'hf0eff43e /* 0x123c */;
            1168: data_o = 32'he575efbf /* 0x1240 */;
            1169: data_o = 32'h00814703 /* 0x1244 */;
            1170: data_o = 32'h04c00793 /* 0x1248 */;
            1171: data_o = 32'h02f71463 /* 0x124c */;
            1172: data_o = 32'h4691480c /* 0x1250 */;
            1173: data_o = 32'h01710713 /* 0x1254 */;
            1174: data_o = 32'h08304785 /* 0x1258 */;
            1175: data_o = 32'hce028522 /* 0x125c */;
            1176: data_o = 32'hd202d002 /* 0x1260 */;
            1177: data_o = 32'hde02dc02 /* 0x1264 */;
            1178: data_o = 32'hf43acc36 /* 0x1268 */;
            1179: data_o = 32'hf0eff83e /* 0x126c */;
            1180: data_o = 32'hed55ecbf /* 0x1270 */;
            1181: data_o = 32'heccef4a6 /* 0x1274 */;
            1182: data_o = 32'h44a1e8d2 /* 0x1278 */;
            1183: data_o = 32'h49854a11 /* 0x127c */;
            1184: data_o = 32'h0783a029 /* 0x1280 */;
            1185: data_o = 32'hdd630009 /* 0x1284 */;
            1186: data_o = 32'h480c0207 /* 0x1288 */;
            1187: data_o = 32'h85220830 /* 0x128c */;
            1188: data_o = 32'hd002ce02 /* 0x1290 */;
            1189: data_o = 32'hdc02d202 /* 0x1294 */;
            1190: data_o = 32'hcc52de02 /* 0x1298 */;
            1191: data_o = 32'hf84ef44a /* 0x129c */;
            1192: data_o = 32'he99ff0ef /* 0x12a0 */;
            1193: data_o = 32'he14934fd /* 0x12a4 */;
            1194: data_o = 32'h74a6fce9 /* 0x12a8 */;
            1195: data_o = 32'h6a4669e6 /* 0x12ac */;
            1196: data_o = 32'h70e64549 /* 0x12b0 */;
            1197: data_o = 32'h79067446 /* 0x12b4 */;
            1198: data_o = 32'h6b066aa6 /* 0x12b8 */;
            1199: data_o = 32'h80826109 /* 0x12bc */;
            1200: data_o = 32'h033b0963 /* 0x12c0 */;
            1201: data_o = 32'h020b1713 /* 0x12c4 */;
            1202: data_o = 32'h01d75b13 /* 0x12c8 */;
            1203: data_o = 32'h16c18793 /* 0x12cc */;
            1204: data_o = 32'h639c97da /* 0x12d0 */;
            1205: data_o = 32'he7b517fd /* 0x12d4 */;
            1206: data_o = 32'h080a8663 /* 0x12d8 */;
            1207: data_o = 32'h744670e6 /* 0x12dc */;
            1208: data_o = 32'h69e674a6 /* 0x12e0 */;
            1209: data_o = 32'h79066a46 /* 0x12e4 */;
            1210: data_o = 32'h6b066aa6 /* 0x12e8 */;
            1211: data_o = 32'h61094501 /* 0x12ec */;
            1212: data_o = 32'h64e18082 /* 0x12f0 */;
            1213: data_o = 32'h6a048493 /* 0x12f4 */;
            1214: data_o = 32'h09934a11 /* 0x12f8 */;
            1215: data_o = 32'h49050171 /* 0x12fc */;
            1216: data_o = 32'hc4ada029 /* 0x1300 */;
            1217: data_o = 32'h01714783 /* 0x1304 */;
            1218: data_o = 32'h480cfbe1 /* 0x1308 */;
            1219: data_o = 32'h85220830 /* 0x130c */;
            1220: data_o = 32'hd002ce02 /* 0x1310 */;
            1221: data_o = 32'hdc02d202 /* 0x1314 */;
            1222: data_o = 32'hcc52de02 /* 0x1318 */;
            1223: data_o = 32'hf84af44e /* 0x131c */;
            1224: data_o = 32'he19ff0ef /* 0x1320 */;
            1225: data_o = 32'hdd7134fd /* 0x1324 */;
            1226: data_o = 32'h69e674a6 /* 0x1328 */;
            1227: data_o = 32'h70e66a46 /* 0x132c */;
            1228: data_o = 32'h79067446 /* 0x1330 */;
            1229: data_o = 32'h6b066aa6 /* 0x1334 */;
            1230: data_o = 32'h6109450d /* 0x1338 */;
            1231: data_o = 32'h46858082 /* 0x133c */;
            1232: data_o = 32'h480cb5d5 /* 0x1340 */;
            1233: data_o = 32'h08300905 /* 0x1344 */;
            1234: data_o = 32'hf44a8522 /* 0x1348 */;
            1235: data_o = 32'hd002ce02 /* 0x134c */;
            1236: data_o = 32'hdc02d202 /* 0x1350 */;
            1237: data_o = 32'hcc52de02 /* 0x1354 */;
            1238: data_o = 32'hf0eff83e /* 0x1358 */;
            1239: data_o = 32'hf569ddff /* 0x135c */;
            1240: data_o = 32'hf60a9ee3 /* 0x1360 */;
            1241: data_o = 32'hf0ef8522 /* 0x1364 */;
            1242: data_o = 32'hbf8dbf7f /* 0x1368 */;
            1243: data_o = 32'h69e674a6 /* 0x136c */;
            1244: data_o = 32'h454d6a46 /* 0x1370 */;
            1245: data_o = 32'h7179bf3d /* 0x1374 */;
            1246: data_o = 32'he84af022 /* 0x1378 */;
            1247: data_o = 32'h8936843a /* 0x137c */;
            1248: data_o = 32'h00344701 /* 0x1380 */;
            1249: data_o = 32'hf406ec26 /* 0x1384 */;
            1250: data_o = 32'hf0ef84b2 /* 0x1388 */;
            1251: data_o = 32'he50de79f /* 0x138c */;
            1252: data_o = 32'h02090463 /* 0x1390 */;
            1253: data_o = 32'h02049713 /* 0x1394 */;
            1254: data_o = 32'h01d75613 /* 0x1398 */;
            1255: data_o = 32'h16c18793 /* 0x139c */;
            1256: data_o = 32'h639897b2 /* 0x13a0 */;
            1257: data_o = 32'h478566a2 /* 0x13a4 */;
            1258: data_o = 32'h0037171b /* 0x13a8 */;
            1259: data_o = 32'h00e797bb /* 0x13ac */;
            1260: data_o = 32'h8c3537fd /* 0x13b0 */;
            1261: data_o = 32'he4198c7d /* 0x13b4 */;
            1262: data_o = 32'h740270a2 /* 0x13b8 */;
            1263: data_o = 32'h694264e2 /* 0x13bc */;
            1264: data_o = 32'h80826145 /* 0x13c0 */;
            1265: data_o = 32'h740270a2 /* 0x13c4 */;
            1266: data_o = 32'h64e28ff5 /* 0x13c8 */;
            1267: data_o = 32'h851b6942 /* 0x13cc */;
            1268: data_o = 32'h61450007 /* 0x13d0 */;
            1269: data_o = 32'h71598082 /* 0x13d4 */;
            1270: data_o = 32'he8caf486 /* 0x13d8 */;
            1271: data_o = 32'h16050963 /* 0x13dc */;
            1272: data_o = 32'h01052903 /* 0x13e0 */;
            1273: data_o = 32'he4cef0a2 /* 0x13e4 */;
            1274: data_o = 32'h842a4989 /* 0x13e8 */;
            1275: data_o = 32'h0729c063 /* 0x13ec */;
            1276: data_o = 32'h016e37b7 /* 0x13f0 */;
            1277: data_o = 32'h8793eca6 /* 0x13f4 */;
            1278: data_o = 32'h84ae5ff7 /* 0x13f8 */;
            1279: data_o = 32'h02b7ff63 /* 0x13fc */;
            1280: data_o = 32'h01003517 /* 0x1400 */;
            1281: data_o = 32'hc0050513 /* 0x1404 */;
            1282: data_o = 32'hf0efe008 /* 0x1408 */;
            1283: data_o = 32'h2481db8f /* 0x140c */;
            1284: data_o = 32'h000315b7 /* 0x1410 */;
            1285: data_o = 32'he002e44a /* 0x1414 */;
            1286: data_o = 32'h85228626 /* 0x1418 */;
            1287: data_o = 32'hd4058593 /* 0x141c */;
            1288: data_o = 32'h48014881 /* 0x1420 */;
            1289: data_o = 32'h47014781 /* 0x1424 */;
            1290: data_o = 32'hf0ef4681 /* 0x1428 */;
            1291: data_o = 32'hc11dd30f /* 0x142c */;
            1292: data_o = 32'h64e67406 /* 0x1430 */;
            1293: data_o = 32'h490d69a6 /* 0x1434 */;
            1294: data_o = 32'h7406a029 /* 0x1438 */;
            1295: data_o = 32'h69a664e6 /* 0x143c */;
            1296: data_o = 32'h70a64961 /* 0x1440 */;
            1297: data_o = 32'h6946854a /* 0x1444 */;
            1298: data_o = 32'h80826165 /* 0x1448 */;
            1299: data_o = 32'h69a67406 /* 0x144c */;
            1300: data_o = 32'hbfc54955 /* 0x1450 */;
            1301: data_o = 32'h15b7485c /* 0x1454 */;
            1302: data_o = 32'he0020003 /* 0x1458 */;
            1303: data_o = 32'h8593e43e /* 0x145c */;
            1304: data_o = 32'h4881d405 /* 0x1460 */;
            1305: data_o = 32'h47814801 /* 0x1464 */;
            1306: data_o = 32'h46814701 /* 0x1468 */;
            1307: data_o = 32'h85228626 /* 0x146c */;
            1308: data_o = 32'hceaff0ef /* 0x1470 */;
            1309: data_o = 32'h3717fd55 /* 0x1474 */;
            1310: data_o = 32'h07130100 /* 0x1478 */;
            1311: data_o = 32'h06b7b8a7 /* 0x147c */;
            1312: data_o = 32'h37978000 /* 0x1480 */;
            1313: data_o = 32'hcb140100 /* 0x1484 */;
            1314: data_o = 32'hb7e78793 /* 0x1488 */;
            1315: data_o = 32'h06b74b98 /* 0x148c */;
            1316: data_o = 32'h37972000 /* 0x1490 */;
            1317: data_o = 32'h87930100 /* 0x1494 */;
            1318: data_o = 32'h8f55b6e7 /* 0x1498 */;
            1319: data_o = 32'h02400613 /* 0x149c */;
            1320: data_o = 32'hcb984581 /* 0x14a0 */;
            1321: data_o = 32'he0ef0868 /* 0x14a4 */;
            1322: data_o = 32'h480ccfff /* 0x14a8 */;
            1323: data_o = 32'h05000793 /* 0x14ac */;
            1324: data_o = 32'h85220830 /* 0x14b0 */;
            1325: data_o = 32'hf43ecc4e /* 0x14b4 */;
            1326: data_o = 32'hc81ff0ef /* 0x14b8 */;
            1327: data_o = 32'h0593f935 /* 0x14bc */;
            1328: data_o = 32'h47050950 /* 0x14c0 */;
            1329: data_o = 32'h859315a2 /* 0x14c4 */;
            1330: data_o = 32'h86ba0405 /* 0x14c8 */;
            1331: data_o = 32'h85224601 /* 0x14cc */;
            1332: data_o = 32'hea7ff0ef /* 0x14d0 */;
            1333: data_o = 32'he925892a /* 0x14d4 */;
            1334: data_o = 32'h0087b5b7 /* 0x14d8 */;
            1335: data_o = 32'ha0158593 /* 0x14dc */;
            1336: data_o = 32'h0aa01737 /* 0x14e0 */;
            1337: data_o = 32'h073205e2 /* 0x14e4 */;
            1338: data_o = 32'h04858593 /* 0x14e8 */;
            1339: data_o = 32'h46850705 /* 0x14ec */;
            1340: data_o = 32'h85224611 /* 0x14f0 */;
            1341: data_o = 32'he83ff0ef /* 0x14f4 */;
            1342: data_o = 32'he531892a /* 0x14f8 */;
            1343: data_o = 32'h07700993 /* 0x14fc */;
            1344: data_o = 32'h098509ea /* 0x1500 */;
            1345: data_o = 32'h478509ba /* 0x1504 */;
            1346: data_o = 32'h06998993 /* 0x1508 */;
            1347: data_o = 32'h00f10c23 /* 0x150c */;
            1348: data_o = 32'hf0efa801 /* 0x1510 */;
            1349: data_o = 32'h892acf1f /* 0x1514 */;
            1350: data_o = 32'h4783e51d /* 0x1518 */;
            1351: data_o = 32'hcb950181 /* 0x151c */;
            1352: data_o = 32'h06500593 /* 0x1520 */;
            1353: data_o = 32'h859315a2 /* 0x1524 */;
            1354: data_o = 32'h47010775 /* 0x1528 */;
            1355: data_o = 32'h46014681 /* 0x152c */;
            1356: data_o = 32'hf0ef8522 /* 0x1530 */;
            1357: data_o = 32'h892ae45f /* 0x1534 */;
            1358: data_o = 32'h08344701 /* 0x1538 */;
            1359: data_o = 32'h85ce4601 /* 0x153c */;
            1360: data_o = 32'h08e38522 /* 0x1540 */;
            1361: data_o = 32'h7406fc09 /* 0x1544 */;
            1362: data_o = 32'h69a664e6 /* 0x1548 */;
            1363: data_o = 32'h4951bddd /* 0x154c */;
            1364: data_o = 32'h0593bdcd /* 0x1550 */;
            1365: data_o = 32'h15a20fd0 /* 0x1554 */;
            1366: data_o = 32'h07a58593 /* 0x1558 */;
            1367: data_o = 32'h46814701 /* 0x155c */;
            1368: data_o = 32'h8522460d /* 0x1560 */;
            1369: data_o = 32'he13ff0ef /* 0x1564 */;
            1370: data_o = 32'hfd71892a /* 0x1568 */;
            1371: data_o = 32'h000a85b7 /* 0x156c */;
            1372: data_o = 32'h05e60585 /* 0x1570 */;
            1373: data_o = 32'h05058593 /* 0x1574 */;
            1374: data_o = 32'h46854701 /* 0x1578 */;
            1375: data_o = 32'h85224601 /* 0x157c */;
            1376: data_o = 32'hf0efe0d2 /* 0x1580 */;
            1377: data_o = 32'h892adf5f /* 0x1584 */;
            1378: data_o = 32'h3983e53d /* 0x1588 */;
            1379: data_o = 32'h07370004 /* 0x158c */;
            1380: data_o = 32'h177de000 /* 0x1590 */;
            1381: data_o = 32'h0109a783 /* 0x1594 */;
            1382: data_o = 32'h00842a03 /* 0x1598 */;
            1383: data_o = 32'h8ff94881 /* 0x159c */;
            1384: data_o = 32'h00f9a823 /* 0x15a0 */;
            1385: data_o = 32'h85d2481c /* 0x15a4 */;
            1386: data_o = 32'he43ee002 /* 0x15a8 */;
            1387: data_o = 32'h47814801 /* 0x15ac */;
            1388: data_o = 32'h46814701 /* 0x15b0 */;
            1389: data_o = 32'h85228626 /* 0x15b4 */;
            1390: data_o = 32'hba2ff0ef /* 0x15b8 */;
            1391: data_o = 32'h485ce91d /* 0x15bc */;
            1392: data_o = 32'he0028626 /* 0x15c0 */;
            1393: data_o = 32'h85d2e43e /* 0x15c4 */;
            1394: data_o = 32'h48818522 /* 0x15c8 */;
            1395: data_o = 32'h47814801 /* 0x15cc */;
            1396: data_o = 32'h46814701 /* 0x15d0 */;
            1397: data_o = 32'hb86ff0ef /* 0x15d4 */;
            1398: data_o = 32'ha783ed09 /* 0x15d8 */;
            1399: data_o = 32'h07370109 /* 0x15dc */;
            1400: data_o = 32'h74062000 /* 0x15e0 */;
            1401: data_o = 32'ha8238fd9 /* 0x15e4 */;
            1402: data_o = 32'h64e600f9 /* 0x15e8 */;
            1403: data_o = 32'h6a0669a6 /* 0x15ec */;
            1404: data_o = 32'h6a06bd89 /* 0x15f0 */;
            1405: data_o = 32'h7406bd35 /* 0x15f4 */;
            1406: data_o = 32'h69a664e6 /* 0x15f8 */;
            1407: data_o = 32'hb5916a06 /* 0x15fc */;
            1408: data_o = 32'hd2010113 /* 0x1600 */;
            1409: data_o = 32'h2b613023 /* 0x1604 */;
            1410: data_o = 32'h00d60b33 /* 0x1608 */;
            1411: data_o = 32'h2c813823 /* 0x160c */;
            1412: data_o = 32'h29713c23 /* 0x1610 */;
            1413: data_o = 32'h29813823 /* 0x1614 */;
            1414: data_o = 32'h2c113c23 /* 0x1618 */;
            1415: data_o = 32'h2c913423 /* 0x161c */;
            1416: data_o = 32'h1ffb7b13 /* 0x1620 */;
            1417: data_o = 32'h8bae842a /* 0x1624 */;
            1418: data_o = 32'h1ff67c13 /* 0x1628 */;
            1419: data_o = 32'h000b1463 /* 0x162c */;
            1420: data_o = 32'h20000b13 /* 0x1630 */;
            1421: data_o = 32'h1ff68493 /* 0x1634 */;
            1422: data_o = 32'h80a594e2 /* 0x1638 */;
            1423: data_o = 32'h34048463 /* 0x163c */;
            1424: data_o = 32'h2d213023 /* 0x1640 */;
            1425: data_o = 32'h8d634785 /* 0x1644 */;
            1426: data_o = 32'h05130cf4 /* 0x1648 */;
            1427: data_o = 32'h82250520 /* 0x164c */;
            1428: data_o = 32'h0ff00693 /* 0x1650 */;
            1429: data_o = 32'h0086579b /* 0x1654 */;
            1430: data_o = 32'h0186559b /* 0x1658 */;
            1431: data_o = 32'h02061713 /* 0x165c */;
            1432: data_o = 32'h8f751682 /* 0x1660 */;
            1433: data_o = 32'h06b707e2 /* 0x1664 */;
            1434: data_o = 32'h05a200ff /* 0x1668 */;
            1435: data_o = 32'h17828e75 /* 0x166c */;
            1436: data_o = 32'h93818dd9 /* 0x1670 */;
            1437: data_o = 32'h8ddd8dd1 /* 0x1674 */;
            1438: data_o = 32'hf8ae8dc9 /* 0x1678 */;
            1439: data_o = 32'h05131894 /* 0x167c */;
            1440: data_o = 32'h47810751 /* 0x1680 */;
            1441: data_o = 32'h0006c603 /* 0x1684 */;
            1442: data_o = 32'h0017979b /* 0x1688 */;
            1443: data_o = 32'hf7938fb1 /* 0x168c */;
            1444: data_o = 32'h87130ff7 /* 0x1690 */;
            1445: data_o = 32'h97ba06c1 /* 0x1694 */;
            1446: data_o = 32'hc7830685 /* 0x1698 */;
            1447: data_o = 32'h93e30007 /* 0x169c */;
            1448: data_o = 32'h979bfea6 /* 0x16a0 */;
            1449: data_o = 32'he7930017 /* 0x16a4 */;
            1450: data_o = 32'h17a20017 /* 0x16a8 */;
            1451: data_o = 32'h04510913 /* 0x16ac */;
            1452: data_o = 32'h86ca8ddd /* 0x16b0 */;
            1453: data_o = 32'h46014705 /* 0x16b4 */;
            1454: data_o = 32'hf0ef8522 /* 0x16b8 */;
            1455: data_o = 32'h1263b49f /* 0x16bc */;
            1456: data_o = 32'h87b31605 /* 0x16c0 */;
            1457: data_o = 32'h3c23418b /* 0x16c4 */;
            1458: data_o = 32'h38232b31 /* 0x16c8 */;
            1459: data_o = 32'h34232b41 /* 0x16cc */;
            1460: data_o = 32'h34232b51 /* 0x16d0 */;
            1461: data_o = 32'h30232991 /* 0x16d4 */;
            1462: data_o = 32'hf43e29a1 /* 0x16d8 */;
            1463: data_o = 32'he402e03e /* 0x16dc */;
            1464: data_o = 32'h4a114c81 /* 0x16e0 */;
            1465: data_o = 32'h0a934985 /* 0x16e4 */;
            1466: data_o = 32'h67e10ff0 /* 0x16e8 */;
            1467: data_o = 32'h6a078d13 /* 0x16ec */;
            1468: data_o = 32'h0a63a039 /* 0x16f0 */;
            1469: data_o = 32'h47031a0d /* 0x16f4 */;
            1470: data_o = 32'h16630451 /* 0x16f8 */;
            1471: data_o = 32'h480c0357 /* 0x16fc */;
            1472: data_o = 32'h852200b0 /* 0x1700 */;
            1473: data_o = 32'hc882c682 /* 0x1704 */;
            1474: data_o = 32'hd482ca82 /* 0x1708 */;
            1475: data_o = 32'hc4d2d682 /* 0x170c */;
            1476: data_o = 32'hf0ceecca /* 0x1710 */;
            1477: data_o = 32'ha25ff0ef /* 0x1714 */;
            1478: data_o = 32'hdd613d7d /* 0x1718 */;
            1479: data_o = 32'ha269450d /* 0x171c */;
            1480: data_o = 32'h05100513 /* 0x1720 */;
            1481: data_o = 32'h0793b72d /* 0x1724 */;
            1482: data_o = 32'h1e630fe0 /* 0x1728 */;
            1483: data_o = 32'h3c2320f7 /* 0x172c */;
            1484: data_o = 32'h896327b1 /* 0x1730 */;
            1485: data_o = 32'h6702100c /* 0x1734 */;
            1486: data_o = 32'hfff48793 /* 0x1738 */;
            1487: data_o = 32'h8063883a /* 0x173c */;
            1488: data_o = 32'h67a21397 /* 0x1740 */;
            1489: data_o = 32'hec02f002 /* 0x1744 */;
            1490: data_o = 32'hf83efc3a /* 0x1748 */;
            1491: data_o = 32'h0d138dc2 /* 0x174c */;
            1492: data_o = 32'h87c22008 /* 0x1750 */;
            1493: data_o = 32'h12078363 /* 0x1754 */;
            1494: data_o = 32'hc4ba4711 /* 0x1758 */;
            1495: data_o = 32'h10000713 /* 0x175c */;
            1496: data_o = 32'hc882c682 /* 0x1760 */;
            1497: data_o = 32'hd482ca82 /* 0x1764 */;
            1498: data_o = 32'hecbed682 /* 0x1768 */;
            1499: data_o = 32'h480cf0ba /* 0x176c */;
            1500: data_o = 32'h852200b0 /* 0x1770 */;
            1501: data_o = 32'hf0efe83e /* 0x1774 */;
            1502: data_o = 32'h67c29c3f /* 0x1778 */;
            1503: data_o = 32'h10078793 /* 0x177c */;
            1504: data_o = 32'h16051c63 /* 0x1780 */;
            1505: data_o = 32'hfda798e3 /* 0x1784 */;
            1506: data_o = 32'h4791480c /* 0x1788 */;
            1507: data_o = 32'h04610713 /* 0x178c */;
            1508: data_o = 32'h00b0c4be /* 0x1790 */;
            1509: data_o = 32'h85224789 /* 0x1794 */;
            1510: data_o = 32'hc882c682 /* 0x1798 */;
            1511: data_o = 32'hd482ca82 /* 0x179c */;
            1512: data_o = 32'hecbad682 /* 0x17a0 */;
            1513: data_o = 32'hf0eff0be /* 0x17a4 */;
            1514: data_o = 32'h1763993f /* 0x17a8 */;
            1515: data_o = 32'h47011405 /* 0x17ac */;
            1516: data_o = 32'h000dc603 /* 0x17b0 */;
            1517: data_o = 32'h0087569b /* 0x17b4 */;
            1518: data_o = 32'h06868eb1 /* 0x17b8 */;
            1519: data_o = 32'he6c18793 /* 0x17bc */;
            1520: data_o = 32'hd78397b6 /* 0x17c0 */;
            1521: data_o = 32'h171b0007 /* 0x17c4 */;
            1522: data_o = 32'h17420087 /* 0x17c8 */;
            1523: data_o = 32'h0d859341 /* 0x17cc */;
            1524: data_o = 32'h9fe38f3d /* 0x17d0 */;
            1525: data_o = 32'h579bfdad /* 0x17d4 */;
            1526: data_o = 32'h171b0087 /* 0x17d8 */;
            1527: data_o = 32'h8fd90087 /* 0x17dc */;
            1528: data_o = 32'h04615703 /* 0x17e0 */;
            1529: data_o = 32'h93c117c2 /* 0x17e4 */;
            1530: data_o = 32'h16f71a63 /* 0x17e8 */;
            1531: data_o = 32'hc7c567e2 /* 0x17ec */;
            1532: data_o = 32'h188c77c2 /* 0x17f0 */;
            1533: data_o = 32'h853395e2 /* 0x17f4 */;
            1534: data_o = 32'h778200fb /* 0x17f8 */;
            1535: data_o = 32'h0633c3ed /* 0x17fc */;
            1536: data_o = 32'he0ef418b /* 0x1800 */;
            1537: data_o = 32'h67829b3f /* 0x1804 */;
            1538: data_o = 32'h87930c85 /* 0x1808 */;
            1539: data_o = 32'he03e2007 /* 0x180c */;
            1540: data_o = 32'h879367a2 /* 0x1810 */;
            1541: data_o = 32'he43e2007 /* 0x1814 */;
            1542: data_o = 32'h0f948b63 /* 0x1818 */;
            1543: data_o = 32'h27813d83 /* 0x181c */;
            1544: data_o = 32'h3903b5e9 /* 0x1820 */;
            1545: data_o = 32'h30832c01 /* 0x1824 */;
            1546: data_o = 32'h34032d81 /* 0x1828 */;
            1547: data_o = 32'h34832d01 /* 0x182c */;
            1548: data_o = 32'h3b032c81 /* 0x1830 */;
            1549: data_o = 32'h3b832a01 /* 0x1834 */;
            1550: data_o = 32'h3c032981 /* 0x1838 */;
            1551: data_o = 32'h01132901 /* 0x183c */;
            1552: data_o = 32'h80822e01 /* 0x1840 */;
            1553: data_o = 32'hee0c09e3 /* 0x1844 */;
            1554: data_o = 32'h0b348263 /* 0x1848 */;
            1555: data_o = 32'hf00277a2 /* 0x184c */;
            1556: data_o = 32'hfc3ef802 /* 0x1850 */;
            1557: data_o = 32'hec3e4785 /* 0x1854 */;
            1558: data_o = 32'h07010813 /* 0x1858 */;
            1559: data_o = 32'h0793bdc5 /* 0x185c */;
            1560: data_o = 32'h0f632000 /* 0x1860 */;
            1561: data_o = 32'hec0208fb /* 0x1864 */;
            1562: data_o = 32'h08136782 /* 0x1868 */;
            1563: data_o = 32'hfc3e0701 /* 0x186c */;
            1564: data_o = 32'hf83e67a2 /* 0x1870 */;
            1565: data_o = 32'hf03e4785 /* 0x1874 */;
            1566: data_o = 32'h6705bdd1 /* 0x1878 */;
            1567: data_o = 32'h80070713 /* 0x187c */;
            1568: data_o = 32'hc6824689 /* 0x1880 */;
            1569: data_o = 32'hca82c882 /* 0x1884 */;
            1570: data_o = 32'hd282d082 /* 0x1888 */;
            1571: data_o = 32'hd682d482 /* 0x188c */;
            1572: data_o = 32'hc4b6ecba /* 0x1890 */;
            1573: data_o = 32'h7782bde9 /* 0x1894 */;
            1574: data_o = 32'h7562d7bd /* 0x1898 */;
            1575: data_o = 32'h188c865a /* 0x189c */;
            1576: data_o = 32'h915fe0ef /* 0x18a0 */;
            1577: data_o = 32'h4565b78d /* 0x18a4 */;
            1578: data_o = 32'h2d813083 /* 0x18a8 */;
            1579: data_o = 32'h2d013403 /* 0x18ac */;
            1580: data_o = 32'h2c013903 /* 0x18b0 */;
            1581: data_o = 32'h2b813983 /* 0x18b4 */;
            1582: data_o = 32'h2b013a03 /* 0x18b8 */;
            1583: data_o = 32'h2a813a83 /* 0x18bc */;
            1584: data_o = 32'h28813c83 /* 0x18c0 */;
            1585: data_o = 32'h28013d03 /* 0x18c4 */;
            1586: data_o = 32'h2c813483 /* 0x18c8 */;
            1587: data_o = 32'h2a013b03 /* 0x18cc */;
            1588: data_o = 32'h29813b83 /* 0x18d0 */;
            1589: data_o = 32'h29013c03 /* 0x18d4 */;
            1590: data_o = 32'h2e010113 /* 0x18d8 */;
            1591: data_o = 32'h06138082 /* 0x18dc */;
            1592: data_o = 32'h06332000 /* 0x18e0 */;
            1593: data_o = 32'he0ef4186 /* 0x18e4 */;
            1594: data_o = 32'hbf318cff /* 0x18e8 */;
            1595: data_o = 32'h20000793 /* 0x18ec */;
            1596: data_o = 32'h04fb0e63 /* 0x18f0 */;
            1597: data_o = 32'hbf8dec26 /* 0x18f4 */;
            1598: data_o = 32'h27813d83 /* 0x18f8 */;
            1599: data_o = 32'hb76d450d /* 0x18fc */;
            1600: data_o = 32'hf0026782 /* 0x1900 */;
            1601: data_o = 32'hfc3eec02 /* 0x1904 */;
            1602: data_o = 32'hf83e67a2 /* 0x1908 */;
            1603: data_o = 32'h4605b581 /* 0x190c */;
            1604: data_o = 32'h04c48963 /* 0x1910 */;
            1605: data_o = 32'h06100593 /* 0x1914 */;
            1606: data_o = 32'h852215a2 /* 0x1918 */;
            1607: data_o = 32'h04c58593 /* 0x191c */;
            1608: data_o = 32'h00b44701 /* 0x1920 */;
            1609: data_o = 32'h8dfff0ef /* 0x1924 */;
            1610: data_o = 32'h2c013903 /* 0x1928 */;
            1611: data_o = 32'h2b813983 /* 0x192c */;
            1612: data_o = 32'h2b013a03 /* 0x1930 */;
            1613: data_o = 32'h2a813a83 /* 0x1934 */;
            1614: data_o = 32'h28813c83 /* 0x1938 */;
            1615: data_o = 32'h28013d03 /* 0x193c */;
            1616: data_o = 32'h27813d83 /* 0x1940 */;
            1617: data_o = 32'h0513b5cd /* 0x1944 */;
            1618: data_o = 32'hbfb90200 /* 0x1948 */;
            1619: data_o = 32'hf00277a2 /* 0x194c */;
            1620: data_o = 32'hfc3ef802 /* 0x1950 */;
            1621: data_o = 32'h0813ec26 /* 0x1954 */;
            1622: data_o = 32'hbbcd0701 /* 0x1958 */;
            1623: data_o = 32'h02100513 /* 0x195c */;
            1624: data_o = 32'h8522b7e1 /* 0x1960 */;
            1625: data_o = 32'hdf8ff0ef /* 0x1964 */;
            1626: data_o = 32'h2c013903 /* 0x1968 */;
            1627: data_o = 32'h2b813983 /* 0x196c */;
            1628: data_o = 32'h2b013a03 /* 0x1970 */;
            1629: data_o = 32'h2a813a83 /* 0x1974 */;
            1630: data_o = 32'h28813c83 /* 0x1978 */;
            1631: data_o = 32'h28013d03 /* 0x197c */;
            1632: data_o = 32'h27813d83 /* 0x1980 */;
            1633: data_o = 32'hb5454501 /* 0x1984 */;
            1634: data_o = 32'hb99dc291 /* 0x1988 */;
            1635: data_o = 32'h80824501 /* 0x198c */;
            1636: data_o = 32'h030007b7 /* 0x1990 */;
            1637: data_o = 32'h87937139 /* 0x1994 */;
            1638: data_o = 32'hf8220007 /* 0x1998 */;
            1639: data_o = 32'h43a4f426 /* 0x199c */;
            1640: data_o = 32'hfc0643e0 /* 0x19a0 */;
            1641: data_o = 32'h14022481 /* 0x19a4 */;
            1642: data_o = 32'h85229001 /* 0x19a8 */;
            1643: data_o = 32'hc8dfe0ef /* 0x19ac */;
            1644: data_o = 32'h85aa4709 /* 0x19b0 */;
            1645: data_o = 32'h04e48b63 /* 0x19b4 */;
            1646: data_o = 32'h8063478d /* 0x19b8 */;
            1647: data_o = 32'h47850af4 /* 0x19bc */;
            1648: data_o = 32'h0af49763 /* 0x19c0 */;
            1649: data_o = 32'h016e37b7 /* 0x19c4 */;
            1650: data_o = 32'h60078793 /* 0x19c8 */;
            1651: data_o = 32'he4020028 /* 0x19cc */;
            1652: data_o = 32'he83ecc02 /* 0x19d0 */;
            1653: data_o = 32'hf0efce3a /* 0x19d4 */;
            1654: data_o = 32'he11da01f /* 0x19d8 */;
            1655: data_o = 32'h3e800513 /* 0x19dc */;
            1656: data_o = 32'h02a40533 /* 0x19e0 */;
            1657: data_o = 32'h000f47b7 /* 0x19e4 */;
            1658: data_o = 32'h24078793 /* 0x19e8 */;
            1659: data_o = 32'h02f55533 /* 0x19ec */;
            1660: data_o = 32'he0ef0505 /* 0x19f0 */;
            1661: data_o = 32'h002c953f /* 0x19f4 */;
            1662: data_o = 32'hd7418513 /* 0x19f8 */;
            1663: data_o = 32'h8c2ff0ef /* 0x19fc */;
            1664: data_o = 32'h744270e2 /* 0x1a00 */;
            1665: data_o = 32'h612174a2 /* 0x1a04 */;
            1666: data_o = 32'h67378082 /* 0x1a08 */;
            1667: data_o = 32'h67b70989 /* 0x1a0c */;
            1668: data_o = 32'he4020262 /* 0x1a10 */;
            1669: data_o = 32'h0713ec02 /* 0x1a14 */;
            1670: data_o = 32'h87937ff7 /* 0x1a18 */;
            1671: data_o = 32'h6463a007 /* 0x1a1c */;
            1672: data_o = 32'h579300a7 /* 0x1a20 */;
            1673: data_o = 32'he83e0025 /* 0x1a24 */;
            1674: data_o = 32'h47850028 /* 0x1a28 */;
            1675: data_o = 32'he0efcc3e /* 0x1a2c */;
            1676: data_o = 32'hf579fb9f /* 0x1a30 */;
            1677: data_o = 32'h15e00793 /* 0x1a34 */;
            1678: data_o = 32'h02f40533 /* 0x1a38 */;
            1679: data_o = 32'h000f47b7 /* 0x1a3c */;
            1680: data_o = 32'h24078793 /* 0x1a40 */;
            1681: data_o = 32'h02f55533 /* 0x1a44 */;
            1682: data_o = 32'he0ef0505 /* 0x1a48 */;
            1683: data_o = 32'h15378fbf /* 0x1a4c */;
            1684: data_o = 32'h002c0200 /* 0x1a50 */;
            1685: data_o = 32'hf7250513 /* 0x1a54 */;
            1686: data_o = 32'h0028b755 /* 0x1a58 */;
            1687: data_o = 32'hf6efe0ef /* 0x1a5c */;
            1688: data_o = 32'h0537f145 /* 0x1a60 */;
            1689: data_o = 32'h002c0200 /* 0x1a64 */;
            1690: data_o = 32'h5ae50513 /* 0x1a68 */;
            1691: data_o = 32'h7442bf41 /* 0x1a6c */;
            1692: data_o = 32'h74a270e2 /* 0x1a70 */;
            1693: data_o = 32'hf06f6121 /* 0x1a74 */;
            1694: data_o = 32'h0000806f /* 0x1a78 */;
            1695: data_o = 32'h00000000 /* 0x1a7c */;
            1696: data_o = 32'h10210000 /* 0x1a80 */;
            1697: data_o = 32'h30632042 /* 0x1a84 */;
            1698: data_o = 32'h50a54084 /* 0x1a88 */;
            1699: data_o = 32'h70e760c6 /* 0x1a8c */;
            1700: data_o = 32'h91298108 /* 0x1a90 */;
            1701: data_o = 32'hb16ba14a /* 0x1a94 */;
            1702: data_o = 32'hd1adc18c /* 0x1a98 */;
            1703: data_o = 32'hf1efe1ce /* 0x1a9c */;
            1704: data_o = 32'h02101231 /* 0x1aa0 */;
            1705: data_o = 32'h22523273 /* 0x1aa4 */;
            1706: data_o = 32'h429452b5 /* 0x1aa8 */;
            1707: data_o = 32'h62d672f7 /* 0x1aac */;
            1708: data_o = 32'h83189339 /* 0x1ab0 */;
            1709: data_o = 32'ha35ab37b /* 0x1ab4 */;
            1710: data_o = 32'hc39cd3bd /* 0x1ab8 */;
            1711: data_o = 32'he3def3ff /* 0x1abc */;
            1712: data_o = 32'h34432462 /* 0x1ac0 */;
            1713: data_o = 32'h14010420 /* 0x1ac4 */;
            1714: data_o = 32'h74c764e6 /* 0x1ac8 */;
            1715: data_o = 32'h548544a4 /* 0x1acc */;
            1716: data_o = 32'hb54ba56a /* 0x1ad0 */;
            1717: data_o = 32'h95098528 /* 0x1ad4 */;
            1718: data_o = 32'hf5cfe5ee /* 0x1ad8 */;
            1719: data_o = 32'hd58dc5ac /* 0x1adc */;
            1720: data_o = 32'h26723653 /* 0x1ae0 */;
            1721: data_o = 32'h06301611 /* 0x1ae4 */;
            1722: data_o = 32'h66f676d7 /* 0x1ae8 */;
            1723: data_o = 32'h46b45695 /* 0x1aec */;
            1724: data_o = 32'ha77ab75b /* 0x1af0 */;
            1725: data_o = 32'h87389719 /* 0x1af4 */;
            1726: data_o = 32'he7fef7df /* 0x1af8 */;
            1727: data_o = 32'hc7bcd79d /* 0x1afc */;
            1728: data_o = 32'h58e548c4 /* 0x1b00 */;
            1729: data_o = 32'h78a76886 /* 0x1b04 */;
            1730: data_o = 32'h18610840 /* 0x1b08 */;
            1731: data_o = 32'h38232802 /* 0x1b0c */;
            1732: data_o = 32'hd9edc9cc /* 0x1b10 */;
            1733: data_o = 32'hf9afe98e /* 0x1b14 */;
            1734: data_o = 32'h99698948 /* 0x1b18 */;
            1735: data_o = 32'hb92ba90a /* 0x1b1c */;
            1736: data_o = 32'h4ad45af5 /* 0x1b20 */;
            1737: data_o = 32'h6a967ab7 /* 0x1b24 */;
            1738: data_o = 32'h0a501a71 /* 0x1b28 */;
            1739: data_o = 32'h2a123a33 /* 0x1b2c */;
            1740: data_o = 32'hcbdcdbfd /* 0x1b30 */;
            1741: data_o = 32'heb9efbbf /* 0x1b34 */;
            1742: data_o = 32'h8b589b79 /* 0x1b38 */;
            1743: data_o = 32'hab1abb3b /* 0x1b3c */;
            1744: data_o = 32'h7c876ca6 /* 0x1b40 */;
            1745: data_o = 32'h5cc54ce4 /* 0x1b44 */;
            1746: data_o = 32'h3c032c22 /* 0x1b48 */;
            1747: data_o = 32'h1c410c60 /* 0x1b4c */;
            1748: data_o = 32'hfd8fedae /* 0x1b50 */;
            1749: data_o = 32'hddcdcdec /* 0x1b54 */;
            1750: data_o = 32'hbd0bad2a /* 0x1b58 */;
            1751: data_o = 32'h9d498d68 /* 0x1b5c */;
            1752: data_o = 32'h6eb67e97 /* 0x1b60 */;
            1753: data_o = 32'h4ef45ed5 /* 0x1b64 */;
            1754: data_o = 32'h2e323e13 /* 0x1b68 */;
            1755: data_o = 32'h0e701e51 /* 0x1b6c */;
            1756: data_o = 32'hefbeff9f /* 0x1b70 */;
            1757: data_o = 32'hcffcdfdd /* 0x1b74 */;
            1758: data_o = 32'haf3abf1b /* 0x1b78 */;
            1759: data_o = 32'h8f789f59 /* 0x1b7c */;
            1760: data_o = 32'h81a99188 /* 0x1b80 */;
            1761: data_o = 32'ha1ebb1ca /* 0x1b84 */;
            1762: data_o = 32'hc12dd10c /* 0x1b88 */;
            1763: data_o = 32'he16ff14e /* 0x1b8c */;
            1764: data_o = 32'h00a11080 /* 0x1b90 */;
            1765: data_o = 32'h20e330c2 /* 0x1b94 */;
            1766: data_o = 32'h40255004 /* 0x1b98 */;
            1767: data_o = 32'h60677046 /* 0x1b9c */;
            1768: data_o = 32'h939883b9 /* 0x1ba0 */;
            1769: data_o = 32'hb3daa3fb /* 0x1ba4 */;
            1770: data_o = 32'hd31cc33d /* 0x1ba8 */;
            1771: data_o = 32'hf35ee37f /* 0x1bac */;
            1772: data_o = 32'h129002b1 /* 0x1bb0 */;
            1773: data_o = 32'h32d222f3 /* 0x1bb4 */;
            1774: data_o = 32'h52144235 /* 0x1bb8 */;
            1775: data_o = 32'h72566277 /* 0x1bbc */;
            1776: data_o = 32'ha5cbb5ea /* 0x1bc0 */;
            1777: data_o = 32'h858995a8 /* 0x1bc4 */;
            1778: data_o = 32'he54ff56e /* 0x1bc8 */;
            1779: data_o = 32'hc50dd52c /* 0x1bcc */;
            1780: data_o = 32'h24c334e2 /* 0x1bd0 */;
            1781: data_o = 32'h048114a0 /* 0x1bd4 */;
            1782: data_o = 32'h64477466 /* 0x1bd8 */;
            1783: data_o = 32'h44055424 /* 0x1bdc */;
            1784: data_o = 32'hb7faa7db /* 0x1be0 */;
            1785: data_o = 32'h97b88799 /* 0x1be4 */;
            1786: data_o = 32'hf77ee75f /* 0x1be8 */;
            1787: data_o = 32'hd73cc71d /* 0x1bec */;
            1788: data_o = 32'h36f226d3 /* 0x1bf0 */;
            1789: data_o = 32'h16b00691 /* 0x1bf4 */;
            1790: data_o = 32'h76766657 /* 0x1bf8 */;
            1791: data_o = 32'h56344615 /* 0x1bfc */;
            1792: data_o = 32'hc96dd94c /* 0x1c00 */;
            1793: data_o = 32'he92ff90e /* 0x1c04 */;
            1794: data_o = 32'h89e999c8 /* 0x1c08 */;
            1795: data_o = 32'ha9abb98a /* 0x1c0c */;
            1796: data_o = 32'h48655844 /* 0x1c10 */;
            1797: data_o = 32'h68277806 /* 0x1c14 */;
            1798: data_o = 32'h08e118c0 /* 0x1c18 */;
            1799: data_o = 32'h28a33882 /* 0x1c1c */;
            1800: data_o = 32'hdb5ccb7d /* 0x1c20 */;
            1801: data_o = 32'hfb1eeb3f /* 0x1c24 */;
            1802: data_o = 32'h9bd88bf9 /* 0x1c28 */;
            1803: data_o = 32'hbb9aabbb /* 0x1c2c */;
            1804: data_o = 32'h5a544a75 /* 0x1c30 */;
            1805: data_o = 32'h7a166a37 /* 0x1c34 */;
            1806: data_o = 32'h1ad00af1 /* 0x1c38 */;
            1807: data_o = 32'h3a922ab3 /* 0x1c3c */;
            1808: data_o = 32'hed0ffd2e /* 0x1c40 */;
            1809: data_o = 32'hcd4ddd6c /* 0x1c44 */;
            1810: data_o = 32'had8bbdaa /* 0x1c48 */;
            1811: data_o = 32'h8dc99de8 /* 0x1c4c */;
            1812: data_o = 32'h6c077c26 /* 0x1c50 */;
            1813: data_o = 32'h4c455c64 /* 0x1c54 */;
            1814: data_o = 32'h2c833ca2 /* 0x1c58 */;
            1815: data_o = 32'h0cc11ce0 /* 0x1c5c */;
            1816: data_o = 32'hff3eef1f /* 0x1c60 */;
            1817: data_o = 32'hdf7ccf5d /* 0x1c64 */;
            1818: data_o = 32'hbfbaaf9b /* 0x1c68 */;
            1819: data_o = 32'h9ff88fd9 /* 0x1c6c */;
            1820: data_o = 32'h7e366e17 /* 0x1c70 */;
            1821: data_o = 32'h5e744e55 /* 0x1c74 */;
            1822: data_o = 32'h3eb22e93 /* 0x1c78 */;
            1823: data_o = 32'h1ef00ed1 /* 0x1c7c */;
            1824: data_o = 32'h36241200 /* 0x1c80 */;
            1825: data_o = 32'h7e6c5a48 /* 0x1c84 */;
            1826: data_o = 32'ha6b48290 /* 0x1c88 */;
            1827: data_o = 32'heefccad8 /* 0x1c8c */;
            1828: data_o = 32'h04162032 /* 0x1c90 */;
            1829: data_o = 32'h4c5e687a /* 0x1c94 */;
            1830: data_o = 32'h9486b0a2 /* 0x1c98 */;
            1831: data_o = 32'hdccef8ea /* 0x1c9c */;
            1832: data_o = 32'h52407664 /* 0x1ca0 */;
            1833: data_o = 32'h1a083e2c /* 0x1ca4 */;
            1834: data_o = 32'hc2d0e6f4 /* 0x1ca8 */;
            1835: data_o = 32'h8a98aebc /* 0x1cac */;
            1836: data_o = 32'h60724456 /* 0x1cb0 */;
            1837: data_o = 32'h283a0c1e /* 0x1cb4 */;
            1838: data_o = 32'hf0e2d4c6 /* 0x1cb8 */;
            1839: data_o = 32'hb8aa9c8e /* 0x1cbc */;
            1840: data_o = 32'hfeecdac8 /* 0x1cc0 */;
            1841: data_o = 32'hb6a49280 /* 0x1cc4 */;
            1842: data_o = 32'h6e7c4a58 /* 0x1cc8 */;
            1843: data_o = 32'h26340210 /* 0x1ccc */;
            1844: data_o = 32'hccdee8fa /* 0x1cd0 */;
            1845: data_o = 32'h8496a0b2 /* 0x1cd4 */;
            1846: data_o = 32'h5c4e786a /* 0x1cd8 */;
            1847: data_o = 32'h14063022 /* 0x1cdc */;
            1848: data_o = 32'h9a88beac /* 0x1ce0 */;
            1849: data_o = 32'hd2c0f6e4 /* 0x1ce4 */;
            1850: data_o = 32'h0a182e3c /* 0x1ce8 */;
            1851: data_o = 32'h42506674 /* 0x1cec */;
            1852: data_o = 32'ha8ba8c9e /* 0x1cf0 */;
            1853: data_o = 32'he0f2c4d6 /* 0x1cf4 */;
            1854: data_o = 32'h382a1c0e /* 0x1cf8 */;
            1855: data_o = 32'h70625446 /* 0x1cfc */;
            1856: data_o = 32'hb4a69082 /* 0x1d00 */;
            1857: data_o = 32'hfceed8ca /* 0x1d04 */;
            1858: data_o = 32'h24360012 /* 0x1d08 */;
            1859: data_o = 32'h6c7e485a /* 0x1d0c */;
            1860: data_o = 32'h8694a2b0 /* 0x1d10 */;
            1861: data_o = 32'hcedceaf8 /* 0x1d14 */;
            1862: data_o = 32'h16043220 /* 0x1d18 */;
            1863: data_o = 32'h5e4c7a68 /* 0x1d1c */;
            1864: data_o = 32'hd0c2f4e6 /* 0x1d20 */;
            1865: data_o = 32'h988abcae /* 0x1d24 */;
            1866: data_o = 32'h40526476 /* 0x1d28 */;
            1867: data_o = 32'h081a2c3e /* 0x1d2c */;
            1868: data_o = 32'he2f0c6d4 /* 0x1d30 */;
            1869: data_o = 32'haab88e9c /* 0x1d34 */;
            1870: data_o = 32'h72605644 /* 0x1d38 */;
            1871: data_o = 32'h3a281e0c /* 0x1d3c */;
            1872: data_o = 32'h7c6e584a /* 0x1d40 */;
            1873: data_o = 32'h34261002 /* 0x1d44 */;
            1874: data_o = 32'hecfec8da /* 0x1d48 */;
            1875: data_o = 32'ha4b68092 /* 0x1d4c */;
            1876: data_o = 32'h4e5c6a78 /* 0x1d50 */;
            1877: data_o = 32'h06142230 /* 0x1d54 */;
            1878: data_o = 32'hdeccfae8 /* 0x1d58 */;
            1879: data_o = 32'h9684b2a0 /* 0x1d5c */;
            1880: data_o = 32'h180a3c2e /* 0x1d60 */;
            1881: data_o = 32'h50427466 /* 0x1d64 */;
            1882: data_o = 32'h889aacbe /* 0x1d68 */;
            1883: data_o = 32'hc0d2e4f6 /* 0x1d6c */;
            1884: data_o = 32'h2a380e1c /* 0x1d70 */;
            1885: data_o = 32'h62704654 /* 0x1d74 */;
            1886: data_o = 32'hbaa89e8c /* 0x1d78 */;
            1887: data_o = 32'hf2e0d6c4 /* 0x1d7c */;
            1888: data_o = 32'h00000001 /* 0x1d80 */;
            1889: data_o = 32'h00000000 /* 0x1d84 */;
            1890: data_o = 32'h00000001 /* 0x1d88 */;
            1891: data_o = 32'h00000000 /* 0x1d8c */;
            1892: data_o = 32'h00000002 /* 0x1d90 */;
            1893: data_o = 32'h00000000 /* 0x1d94 */;
            1894: data_o = 32'h00000005 /* 0x1d98 */;
            1895: data_o = 32'h00000000 /* 0x1d9c */;
            1896: data_o = 32'h00000005 /* 0x1da0 */;
            1897: data_o = 32'h00000000 /* 0x1da4 */;
            1898: data_o = 32'h00000000 /* 0x1da8 */;
            1899: data_o = 32'h00000000 /* 0x1dac */;
            1900: data_o = 32'h00000000 /* 0x1db0 */;
            1901: data_o = 32'h00000000 /* 0x1db4 */;
            1902: data_o = 32'h00000000 /* 0x1db8 */;
            1903: data_o = 32'h00000000 /* 0x1dbc */;
            1904: data_o = 32'h00000000 /* 0x1dc0 */;
            1905: data_o = 32'h00000000 /* 0x1dc4 */;
            1906: data_o = 32'h00000000 /* 0x1dc8 */;
            1907: data_o = 32'h00000000 /* 0x1dcc */;
            1908: data_o = 32'h00000000 /* 0x1dd0 */;
            1909: data_o = 32'h00000000 /* 0x1dd4 */;
            1910: data_o = 32'h00000000 /* 0x1dd8 */;
            1911: data_o = 32'h00000000 /* 0x1ddc */;
            1912: data_o = 32'h00000000 /* 0x1de0 */;
            1913: data_o = 32'h00000000 /* 0x1de4 */;
            1914: data_o = 32'h00000000 /* 0x1de8 */;
            1915: data_o = 32'h00000000 /* 0x1dec */;
            1916: data_o = 32'h00000000 /* 0x1df0 */;
            1917: data_o = 32'h00000000 /* 0x1df4 */;
            1918: data_o = 32'h00000000 /* 0x1df8 */;
            1919: data_o = 32'h00000000 /* 0x1dfc */;
            1920: data_o = 32'h00000000 /* 0x1e00 */;
            1921: data_o = 32'h00000000 /* 0x1e04 */;
            1922: data_o = 32'h00000000 /* 0x1e08 */;
            1923: data_o = 32'h00000000 /* 0x1e0c */;
            1924: data_o = 32'h00000000 /* 0x1e10 */;
            1925: data_o = 32'h00000000 /* 0x1e14 */;
            1926: data_o = 32'h00000000 /* 0x1e18 */;
            1927: data_o = 32'h00000000 /* 0x1e1c */;
            1928: data_o = 32'h00000000 /* 0x1e20 */;
            1929: data_o = 32'h00000000 /* 0x1e24 */;
            1930: data_o = 32'h00000000 /* 0x1e28 */;
            1931: data_o = 32'h00000000 /* 0x1e2c */;
            1932: data_o = 32'h00000000 /* 0x1e30 */;
            1933: data_o = 32'h00000000 /* 0x1e34 */;
            1934: data_o = 32'h00000000 /* 0x1e38 */;
            1935: data_o = 32'h00000000 /* 0x1e3c */;
            1936: data_o = 32'h00000000 /* 0x1e40 */;
            1937: data_o = 32'h00000000 /* 0x1e44 */;
            1938: data_o = 32'h00000000 /* 0x1e48 */;
            1939: data_o = 32'h00000000 /* 0x1e4c */;
            1940: data_o = 32'h00000000 /* 0x1e50 */;
            1941: data_o = 32'h00000000 /* 0x1e54 */;
            1942: data_o = 32'h00000000 /* 0x1e58 */;
            1943: data_o = 32'h00000000 /* 0x1e5c */;
            1944: data_o = 32'h00000000 /* 0x1e60 */;
            1945: data_o = 32'h00000000 /* 0x1e64 */;
            1946: data_o = 32'h00000000 /* 0x1e68 */;
            1947: data_o = 32'h00000000 /* 0x1e6c */;
            1948: data_o = 32'h00000000 /* 0x1e70 */;
            1949: data_o = 32'h00000000 /* 0x1e74 */;
            1950: data_o = 32'h00000000 /* 0x1e78 */;
            1951: data_o = 32'h00000000 /* 0x1e7c */;
            1952: data_o = 32'h00000000 /* 0x1e80 */;
            1953: data_o = 32'h00000000 /* 0x1e84 */;
            1954: data_o = 32'h00000000 /* 0x1e88 */;
            1955: data_o = 32'h00000000 /* 0x1e8c */;
            1956: data_o = 32'h00000000 /* 0x1e90 */;
            1957: data_o = 32'h00000000 /* 0x1e94 */;
            1958: data_o = 32'h00000000 /* 0x1e98 */;
            1959: data_o = 32'h00000000 /* 0x1e9c */;
            1960: data_o = 32'h00000000 /* 0x1ea0 */;
            1961: data_o = 32'h00000000 /* 0x1ea4 */;
            1962: data_o = 32'h00000000 /* 0x1ea8 */;
            1963: data_o = 32'h00000000 /* 0x1eac */;
            1964: data_o = 32'h00000000 /* 0x1eb0 */;
            1965: data_o = 32'h00000000 /* 0x1eb4 */;
            1966: data_o = 32'h00000000 /* 0x1eb8 */;
            1967: data_o = 32'h00000000 /* 0x1ebc */;
            1968: data_o = 32'h00000000 /* 0x1ec0 */;
            1969: data_o = 32'h00000000 /* 0x1ec4 */;
            1970: data_o = 32'h00000000 /* 0x1ec8 */;
            1971: data_o = 32'h00000000 /* 0x1ecc */;
            1972: data_o = 32'h00000000 /* 0x1ed0 */;
            1973: data_o = 32'h00000000 /* 0x1ed4 */;
            1974: data_o = 32'h00000000 /* 0x1ed8 */;
            1975: data_o = 32'h00000000 /* 0x1edc */;
            1976: data_o = 32'h00000000 /* 0x1ee0 */;
            1977: data_o = 32'h00000000 /* 0x1ee4 */;
            1978: data_o = 32'h00000000 /* 0x1ee8 */;
            1979: data_o = 32'h00000000 /* 0x1eec */;
            1980: data_o = 32'h00000000 /* 0x1ef0 */;
            1981: data_o = 32'h00000000 /* 0x1ef4 */;
            1982: data_o = 32'h00000000 /* 0x1ef8 */;
            1983: data_o = 32'h00000000 /* 0x1efc */;
            1984: data_o = 32'h00000000 /* 0x1f00 */;
            1985: data_o = 32'h00000000 /* 0x1f04 */;
            1986: data_o = 32'h00000000 /* 0x1f08 */;
            1987: data_o = 32'h00000000 /* 0x1f0c */;
            1988: data_o = 32'h00000000 /* 0x1f10 */;
            1989: data_o = 32'h00000000 /* 0x1f14 */;
            1990: data_o = 32'h00000000 /* 0x1f18 */;
            1991: data_o = 32'h00000000 /* 0x1f1c */;
            1992: data_o = 32'h00000000 /* 0x1f20 */;
            1993: data_o = 32'h00000000 /* 0x1f24 */;
            1994: data_o = 32'h00000000 /* 0x1f28 */;
            1995: data_o = 32'h00000000 /* 0x1f2c */;
            1996: data_o = 32'h00000000 /* 0x1f30 */;
            1997: data_o = 32'h00000000 /* 0x1f34 */;
            1998: data_o = 32'h00000000 /* 0x1f38 */;
            1999: data_o = 32'h00000000 /* 0x1f3c */;
            2000: data_o = 32'h00000000 /* 0x1f40 */;
            2001: data_o = 32'h00000000 /* 0x1f44 */;
            2002: data_o = 32'h00000000 /* 0x1f48 */;
            2003: data_o = 32'h00000000 /* 0x1f4c */;
            2004: data_o = 32'h00000000 /* 0x1f50 */;
            2005: data_o = 32'h00000000 /* 0x1f54 */;
            2006: data_o = 32'h00000000 /* 0x1f58 */;
            2007: data_o = 32'h00000000 /* 0x1f5c */;
            2008: data_o = 32'h00000000 /* 0x1f60 */;
            2009: data_o = 32'h00000000 /* 0x1f64 */;
            2010: data_o = 32'h00000000 /* 0x1f68 */;
            2011: data_o = 32'h00000000 /* 0x1f6c */;
            2012: data_o = 32'h00000000 /* 0x1f70 */;
            2013: data_o = 32'h00000000 /* 0x1f74 */;
            2014: data_o = 32'h00000000 /* 0x1f78 */;
            2015: data_o = 32'h00000000 /* 0x1f7c */;
            2016: data_o = 32'h00000000 /* 0x1f80 */;
            2017: data_o = 32'h00000000 /* 0x1f84 */;
            2018: data_o = 32'h00000000 /* 0x1f88 */;
            2019: data_o = 32'h00000000 /* 0x1f8c */;
            2020: data_o = 32'h00000000 /* 0x1f90 */;
            2021: data_o = 32'h00000000 /* 0x1f94 */;
            2022: data_o = 32'h00000000 /* 0x1f98 */;
            2023: data_o = 32'h00000000 /* 0x1f9c */;
            2024: data_o = 32'h00000000 /* 0x1fa0 */;
            2025: data_o = 32'h00000000 /* 0x1fa4 */;
            2026: data_o = 32'h00000000 /* 0x1fa8 */;
            2027: data_o = 32'h00000000 /* 0x1fac */;
            2028: data_o = 32'h00000000 /* 0x1fb0 */;
            2029: data_o = 32'h00000000 /* 0x1fb4 */;
            2030: data_o = 32'h00000000 /* 0x1fb8 */;
            2031: data_o = 32'h00000000 /* 0x1fbc */;
            2032: data_o = 32'h00000000 /* 0x1fc0 */;
            2033: data_o = 32'h00000000 /* 0x1fc4 */;
            2034: data_o = 32'h00000000 /* 0x1fc8 */;
            2035: data_o = 32'h00000000 /* 0x1fcc */;
            2036: data_o = 32'h00000000 /* 0x1fd0 */;
            2037: data_o = 32'h00000000 /* 0x1fd4 */;
            2038: data_o = 32'h00000000 /* 0x1fd8 */;
            2039: data_o = 32'h00000000 /* 0x1fdc */;
            2040: data_o = 32'h00000000 /* 0x1fe0 */;
            2041: data_o = 32'h00000000 /* 0x1fe4 */;
            2042: data_o = 32'h00000000 /* 0x1fe8 */;
            2043: data_o = 32'h00000000 /* 0x1fec */;
            2044: data_o = 32'h00000000 /* 0x1ff0 */;
            2045: data_o = 32'h00000000 /* 0x1ff4 */;
            2046: data_o = 32'h00000000 /* 0x1ff8 */;
            2047: data_o = 32'h00000000 /* 0x1ffc */;
            default: data_o = '0;
        endcase
    end

endmodule
